library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ram is port(
    clk   : in  std_logic;
    wr    : in  std_logic;
    addr  : in  std_logic_vector(14 downto 0);
    din   : in  std_logic_vector( 7 downto 0);
    dout  : out std_logic_vector( 7 downto 0));
end ram;

architecture behavioral of ram is

  type ram_t is array (0 to 32767) of std_logic_vector(7 downto 0);
  signal ram : ram_t := (
  X"F3", X"01", X"2B", X"69", X"0B", X"78", X"B1", X"20", --0000
  X"FB", X"C3", X"C7", X"00", X"00", X"00", X"00", X"00", --0008
  X"EF", X"10", X"00", X"C9", X"00", X"00", X"00", X"00", --0010
  X"EF", X"18", X"00", X"C9", X"00", X"00", X"00", X"00", --0018
  X"EF", X"20", X"00", X"C9", X"00", X"00", X"00", X"00", --0020
  X"E3", X"F5", X"7E", X"23", X"23", X"22", X"5A", X"5B", --0028
  X"2B", X"66", X"6F", X"F1", X"C3", X"5C", X"00", X"00", --0030
  X"E5", X"21", X"48", X"00", X"E5", X"21", X"00", X"5B", --0038
  X"E5", X"21", X"38", X"00", X"E5", X"C3", X"00", X"5B", --0040
  X"E1", X"C9", X"01", X"FD", X"7F", X"AF", X"F3", X"ED", --0048
  X"79", X"32", X"5C", X"5B", X"FB", X"3D", X"FD", X"77", --0050
  X"00", X"C3", X"21", X"03", X"22", X"58", X"5B", X"21", --0058
  X"14", X"5B", X"E3", X"E5", X"2A", X"58", X"5B", X"E3", --0060
  X"C3", X"00", X"5B", X"F5", X"C5", X"01", X"FD", X"7F", --0068
  X"3A", X"5C", X"5B", X"EE", X"10", X"F3", X"32", X"5C", --0070
  X"5B", X"ED", X"79", X"FB", X"C1", X"F1", X"C9", X"CD", --0078
  X"00", X"5B", X"E5", X"2A", X"5A", X"5B", X"E3", X"C9", --0080
  X"F3", X"3A", X"5C", X"5B", X"E6", X"EF", X"32", X"5C", --0088
  X"5B", X"01", X"FD", X"7F", X"ED", X"79", X"FB", X"C3", --0090
  X"C3", X"00", X"21", X"D8", X"06", X"18", X"03", X"21", --0098
  X"CA", X"07", X"08", X"01", X"FD", X"7F", X"3A", X"5C", --00A0
  X"5B", X"F5", X"E6", X"EF", X"F3", X"32", X"5C", X"5B", --00A8
  X"ED", X"79", X"C3", X"E6", X"05", X"08", X"F1", X"01", --00B0
  X"FD", X"7F", X"F3", X"32", X"5C", X"5B", X"ED", X"79", --00B8
  X"FB", X"08", X"C9", X"2A", X"8B", X"5B", X"E9", X"06", --00C0
  X"08", X"78", X"D9", X"3D", X"01", X"FD", X"7F", X"ED", --00C8
  X"79", X"21", X"00", X"C0", X"11", X"01", X"C0", X"01", --00D0
  X"FF", X"3F", X"3E", X"FF", X"77", X"BE", X"20", X"51", --00D8
  X"AF", X"77", X"BE", X"20", X"4C", X"ED", X"B0", X"D9", --00E0
  X"10", X"DF", X"32", X"88", X"5B", X"0E", X"FD", X"16", --00E8
  X"FF", X"1E", X"BF", X"42", X"3E", X"0E", X"ED", X"79", --00F0
  X"43", X"3E", X"FF", X"ED", X"79", X"18", X"38", X"00", --00F8
  X"C3", X"AF", X"17", X"C3", X"38", X"18", X"C3", X"CF", --0100
  X"1E", X"C3", X"04", X"1F", X"C3", X"4A", X"00", X"C3", --0108
  X"A2", X"03", X"C3", X"2A", X"18", X"C3", X"A8", X"18", --0110
  X"C3", X"2D", X"01", X"C3", X"05", X"0A", X"C3", X"A3", --0118
  X"11", X"C3", X"D8", X"06", X"C3", X"CA", X"07", X"C3", --0120
  X"A3", X"08", X"C3", X"F0", X"08", X"EF", X"01", X"3B", --0128
  X"C9", X"D9", X"78", X"D3", X"FE", X"18", X"FE", X"42", --0130
  X"3E", X"07", X"ED", X"79", X"43", X"3E", X"FF", X"ED", --0138
  X"79", X"11", X"00", X"5B", X"21", X"6B", X"00", X"01", --0140
  X"58", X"00", X"ED", X"B0", X"3E", X"CF", X"32", X"5D", --0148
  X"5B", X"31", X"FF", X"5B", X"3E", X"04", X"CD", X"64", --0150
  X"1C", X"DD", X"21", X"EC", X"EB", X"DD", X"22", X"83", --0158
  X"5B", X"DD", X"36", X"0A", X"00", X"DD", X"36", X"0B", --0160
  X"C0", X"DD", X"36", X"0C", X"00", X"21", X"EC", X"2B", --0168
  X"3E", X"01", X"22", X"85", X"5B", X"32", X"87", X"5B", --0170
  X"3E", X"05", X"CD", X"64", X"1C", X"21", X"FF", X"FF", --0178
  X"22", X"B4", X"5C", X"11", X"AF", X"3E", X"01", X"A8", --0180
  X"00", X"EB", X"EF", X"61", X"16", X"EB", X"23", X"22", --0188
  X"7B", X"5C", X"2B", X"01", X"40", X"00", X"ED", X"43", --0190
  X"38", X"5C", X"22", X"B2", X"5C", X"21", X"00", X"3C", --0198
  X"22", X"36", X"5C", X"2A", X"B2", X"5C", X"23", X"F9", --01A0
  X"ED", X"56", X"FD", X"21", X"3A", X"5C", X"FD", X"CB", --01A8
  X"01", X"E6", X"FB", X"21", X"0B", X"00", X"22", X"5F", --01B0
  X"5B", X"AF", X"32", X"61", X"5B", X"32", X"63", X"5B", --01B8
  X"32", X"65", X"5B", X"21", X"00", X"EC", X"22", X"24", --01C0
  X"FF", X"3E", X"50", X"32", X"64", X"5B", X"21", X"0A", --01C8
  X"00", X"22", X"94", X"5B", X"22", X"96", X"5B", X"21", --01D0
  X"B6", X"5C", X"22", X"4F", X"5C", X"11", X"89", X"05", --01D8
  X"01", X"15", X"00", X"EB", X"ED", X"B0", X"EB", X"2B", --01E0
  X"22", X"57", X"5C", X"23", X"22", X"53", X"5C", X"22", --01E8
  X"4B", X"5C", X"36", X"80", X"23", X"22", X"59", X"5C", --01F0
  X"36", X"0D", X"23", X"36", X"80", X"23", X"22", X"61", --01F8
  X"5C", X"22", X"63", X"5C", X"22", X"65", X"5C", X"3E", --0200
  X"38", X"32", X"8D", X"5C", X"32", X"8F", X"5C", X"32", --0208
  X"48", X"5C", X"AF", X"32", X"13", X"EC", X"3E", X"07", --0210
  X"D3", X"FE", X"21", X"23", X"05", X"22", X"09", X"5C", --0218
  X"FD", X"35", X"C6", X"FD", X"35", X"CA", X"21", X"9E", --0220
  X"05", X"11", X"10", X"5C", X"01", X"0E", X"00", X"ED", --0228
  X"B0", X"FD", X"CB", X"01", X"8E", X"FD", X"36", X"00", --0230
  X"FF", X"FD", X"36", X"31", X"02", X"EF", X"6B", X"0D", --0238
  X"EF", X"04", X"3C", X"11", X"61", X"05", X"CD", X"7D", --0240
  X"05", X"FD", X"36", X"31", X"02", X"FD", X"CB", X"02", --0248
  X"EE", X"21", X"FF", X"5B", X"22", X"81", X"5B", X"CD", --0250
  X"45", X"1F", X"3E", X"38", X"32", X"11", X"EC", X"32", --0258
  X"0F", X"EC", X"CD", X"84", X"25", X"CD", X"20", X"1F", --0260
  X"C3", X"9F", X"25", X"21", X"66", X"5B", X"CB", X"C6", --0268
  X"FD", X"36", X"00", X"FF", X"FD", X"36", X"31", X"02", --0270
  X"21", X"1D", X"5B", X"E5", X"ED", X"73", X"3D", X"5C", --0278
  X"21", X"BA", X"02", X"22", X"8B", X"5B", X"CD", X"8E", --0280
  X"22", X"CD", X"CB", X"22", X"CA", X"F8", X"21", X"FE", --0288
  X"28", X"CA", X"F8", X"21", X"FE", X"2D", X"CA", X"F8", --0290
  X"21", X"FE", X"2B", X"CA", X"F8", X"21", X"CD", X"E0", --0298
  X"22", X"CA", X"F8", X"21", X"CD", X"45", X"1F", X"3A", --02A0
  X"0E", X"EC", X"CD", X"20", X"1F", X"FE", X"04", X"C2", --02A8
  X"AF", X"17", X"CD", X"97", X"22", X"CA", X"AF", X"17", --02B0
  X"E1", X"C9", X"FD", X"CB", X"00", X"7E", X"20", X"01", --02B8
  X"C9", X"2A", X"59", X"5C", X"22", X"5D", X"5C", X"EF", --02C0
  X"FB", X"19", X"78", X"B1", X"C2", X"F7", X"03", X"DF", --02C8
  X"FE", X"0D", X"C8", X"CD", X"EF", X"21", X"FD", X"CB", --02D0
  X"02", X"76", X"20", X"03", X"EF", X"6E", X"0D", X"FD", --02D8
  X"CB", X"02", X"B6", X"CD", X"45", X"1F", X"21", X"0D", --02E0
  X"EC", X"CB", X"76", X"20", X"07", X"23", X"7E", X"FE", --02E8
  X"00", X"CC", X"81", X"38", X"CD", X"20", X"1F", X"21", --02F0
  X"3C", X"5C", X"CB", X"9E", X"3E", X"19", X"FD", X"96", --02F8
  X"4F", X"32", X"8C", X"5C", X"FD", X"CB", X"01", X"FE", --0300
  X"FD", X"36", X"0A", X"01", X"21", X"00", X"3E", X"E5", --0308
  X"21", X"1D", X"5B", X"E5", X"ED", X"73", X"3D", X"5C", --0310
  X"21", X"21", X"03", X"22", X"8B", X"5B", X"C3", X"38", --0318
  X"18", X"ED", X"7B", X"B2", X"5C", X"33", X"21", X"FF", --0320
  X"5B", X"22", X"81", X"5B", X"76", X"FD", X"CB", X"01", --0328
  X"AE", X"21", X"66", X"5B", X"CB", X"56", X"28", X"12", --0330
  X"CD", X"45", X"1F", X"DD", X"2A", X"83", X"5B", X"01", --0338
  X"14", X"00", X"DD", X"09", X"CD", X"56", X"1D", X"CD", --0340
  X"20", X"1F", X"3A", X"3A", X"5C", X"3C", X"F5", X"21", --0348
  X"00", X"00", X"FD", X"74", X"37", X"FD", X"74", X"26", --0350
  X"22", X"0B", X"5C", X"21", X"01", X"00", X"22", X"16", --0358
  X"5C", X"EF", X"B0", X"16", X"FD", X"CB", X"37", X"AE", --0360
  X"EF", X"6E", X"0D", X"FD", X"CB", X"02", X"EE", X"F1", --0368
  X"47", X"FE", X"0A", X"38", X"0A", X"FE", X"1D", X"38", --0370
  X"04", X"C6", X"14", X"18", X"02", X"C6", X"07", X"EF", --0378
  X"EF", X"15", X"3E", X"20", X"D7", X"78", X"FE", X"1D", --0380
  X"38", X"12", X"D6", X"1D", X"06", X"00", X"4F", X"21", --0388
  X"6C", X"04", X"09", X"09", X"5E", X"23", X"56", X"CD", --0390
  X"7D", X"05", X"18", X"06", X"11", X"91", X"13", X"EF", --0398
  X"0A", X"0C", X"AF", X"11", X"36", X"15", X"EF", X"0A", --03A0
  X"0C", X"ED", X"4B", X"45", X"5C", X"EF", X"1B", X"1A", --03A8
  X"3E", X"3A", X"D7", X"FD", X"4E", X"0D", X"06", X"00", --03B0
  X"EF", X"1B", X"1A", X"EF", X"97", X"10", X"3A", X"3A", --03B8
  X"5C", X"3C", X"28", X"1B", X"FE", X"09", X"28", X"04", --03C0
  X"FE", X"15", X"20", X"03", X"FD", X"34", X"0D", X"01", --03C8
  X"03", X"00", X"11", X"70", X"5C", X"21", X"44", X"5C", --03D0
  X"CB", X"7E", X"28", X"01", X"09", X"ED", X"B8", X"FD", --03D8
  X"36", X"0A", X"FF", X"FD", X"CB", X"01", X"9E", X"21", --03E0
  X"66", X"5B", X"CB", X"86", X"C3", X"CB", X"25", X"3E", --03E8
  X"10", X"01", X"00", X"00", X"C3", X"4E", X"03", X"ED", --03F0
  X"43", X"49", X"5C", X"CD", X"45", X"1F", X"78", X"B1", --03F8
  X"28", X"08", X"ED", X"43", X"49", X"5C", X"ED", X"43", --0400
  X"08", X"EC", X"CD", X"20", X"1F", X"2A", X"5D", X"5C", --0408
  X"EB", X"21", X"EF", X"03", X"E5", X"2A", X"61", X"5C", --0410
  X"37", X"ED", X"52", X"E5", X"60", X"69", X"EF", X"6E", --0418
  X"19", X"20", X"06", X"EF", X"B8", X"19", X"EF", X"E8", --0420
  X"19", X"C1", X"79", X"3D", X"B0", X"20", X"13", X"CD", --0428
  X"45", X"1F", X"E5", X"2A", X"49", X"5C", X"CD", X"4A", --0430
  X"33", X"22", X"49", X"5C", X"E1", X"CD", X"20", X"1F", --0438
  X"18", X"28", X"C5", X"03", X"03", X"03", X"03", X"2B", --0440
  X"ED", X"5B", X"53", X"5C", X"D5", X"EF", X"55", X"16", --0448
  X"E1", X"22", X"53", X"5C", X"C1", X"C5", X"13", X"2A", --0450
  X"61", X"5C", X"2B", X"2B", X"ED", X"B8", X"2A", X"49", --0458
  X"5C", X"EB", X"C1", X"70", X"2B", X"71", X"2B", X"73", --0460
  X"2B", X"72", X"F1", X"C9", X"8C", X"04", X"97", X"04", --0468
  X"A6", X"04", X"B0", X"04", X"C1", X"04", X"D4", X"04", --0470
  X"E0", X"04", X"E0", X"04", X"F3", X"04", X"01", X"05", --0478
  X"12", X"05", X"23", X"05", X"31", X"05", X"42", X"05", --0480
  X"4E", X"05", X"61", X"05", X"4D", X"45", X"52", X"47", --0488
  X"45", X"20", X"65", X"72", X"72", X"6F", X"F2", X"57", --0490
  X"72", X"6F", X"6E", X"67", X"20", X"66", X"69", X"6C", --0498
  X"65", X"20", X"74", X"79", X"70", X"E5", X"43", X"4F", --04A0
  X"44", X"45", X"20", X"65", X"72", X"72", X"6F", X"F2", --04A8
  X"54", X"6F", X"6F", X"20", X"6D", X"61", X"6E", X"79", --04B0
  X"20", X"62", X"72", X"61", X"63", X"6B", X"65", X"74", --04B8
  X"F3", X"46", X"69", X"6C", X"65", X"20", X"61", X"6C", --04C0
  X"72", X"65", X"61", X"64", X"79", X"20", X"65", X"78", --04C8
  X"69", X"73", X"74", X"F3", X"49", X"6E", X"76", X"61", --04D0
  X"6C", X"69", X"64", X"20", X"6E", X"61", X"6D", X"E5", --04D8
  X"46", X"69", X"6C", X"65", X"20", X"64", X"6F", X"65", --04E0
  X"73", X"20", X"6E", X"6F", X"74", X"20", X"65", X"78", --04E8
  X"69", X"73", X"F4", X"49", X"6E", X"76", X"61", X"6C", --04F0
  X"69", X"64", X"20", X"64", X"65", X"76", X"69", X"63", --04F8
  X"E5", X"49", X"6E", X"76", X"61", X"6C", X"69", X"64", --0500
  X"20", X"62", X"61", X"75", X"64", X"20", X"72", X"61", --0508
  X"74", X"E5", X"49", X"6E", X"76", X"61", X"6C", X"69", --0510
  X"64", X"20", X"6E", X"6F", X"74", X"65", X"20", X"6E", --0518
  X"61", X"6D", X"E5", X"4E", X"75", X"6D", X"62", X"65", --0520
  X"72", X"20", X"74", X"6F", X"6F", X"20", X"62", X"69", --0528
  X"E7", X"4E", X"6F", X"74", X"65", X"20", X"6F", X"75", --0530
  X"74", X"20", X"6F", X"66", X"20", X"72", X"61", X"6E", --0538
  X"67", X"E5", X"4F", X"75", X"74", X"20", X"6F", X"66", --0540
  X"20", X"72", X"61", X"6E", X"67", X"E5", X"54", X"6F", --0548
  X"6F", X"20", X"6D", X"61", X"6E", X"79", X"20", X"74", --0550
  X"69", X"65", X"64", X"20", X"6E", X"6F", X"74", X"65", --0558
  X"F3", X"7F", X"20", X"31", X"39", X"38", X"36", X"20", --0560
  X"53", X"69", X"6E", X"63", X"6C", X"61", X"69", X"72", --0568
  X"20", X"52", X"65", X"73", X"65", X"61", X"72", X"63", --0570
  X"68", X"20", X"4C", X"74", X"E4", X"1A", X"E6", X"7F", --0578
  X"D5", X"D7", X"D1", X"1A", X"13", X"87", X"30", X"F5", --0580
  X"C9", X"F4", X"09", X"A8", X"10", X"4B", X"F4", X"09", --0588
  X"C4", X"15", X"53", X"81", X"0F", X"C4", X"15", X"52", --0590
  X"34", X"5B", X"2F", X"5B", X"50", X"80", X"01", X"00", --0598
  X"06", X"00", X"0B", X"00", X"01", X"00", X"01", X"00", --05A0
  X"06", X"00", X"10", X"00", X"E1", X"01", X"FD", X"7F", --05A8
  X"AF", X"F3", X"32", X"5C", X"5B", X"ED", X"79", X"FB", --05B0
  X"ED", X"7B", X"3D", X"5C", X"7E", X"32", X"5E", X"5B", --05B8
  X"3C", X"FE", X"1E", X"30", X"03", X"EF", X"5D", X"5B", --05C0
  X"3D", X"FD", X"77", X"00", X"2A", X"5D", X"5C", X"22", --05C8
  X"5F", X"5C", X"EF", X"C5", X"16", X"C9", X"3E", X"7F", --05D0
  X"DB", X"FE", X"1F", X"D8", X"3E", X"FE", X"DB", X"FE", --05D8
  X"1F", X"D8", X"CD", X"AC", X"05", X"14", X"FB", X"08", --05E0
  X"11", X"4A", X"5B", X"D5", X"FD", X"CB", X"02", X"9E", --05E8
  X"E5", X"2A", X"3D", X"5C", X"5E", X"23", X"56", X"A7", --05F0
  X"21", X"7F", X"10", X"ED", X"52", X"20", X"38", X"E1", --05F8
  X"ED", X"7B", X"3D", X"5C", X"D1", X"D1", X"ED", X"53", --0600
  X"3D", X"5C", X"E5", X"11", X"10", X"06", X"D5", X"E9", --0608
  X"38", X"09", X"28", X"04", X"CD", X"AC", X"05", X"07", --0610
  X"E1", X"18", X"EF", X"FE", X"0D", X"28", X"0E", X"2A", --0618
  X"5A", X"5B", X"E5", X"EF", X"85", X"0F", X"E1", X"22", --0620
  X"5A", X"5B", X"E1", X"18", X"DD", X"E1", X"3A", X"5C", --0628
  X"5B", X"F6", X"10", X"F5", X"C3", X"4A", X"5B", X"E1", --0630
  X"11", X"3D", X"06", X"D5", X"E9", X"D8", X"C8", X"18", --0638
  X"D3", X"EF", X"18", X"00", X"EF", X"8C", X"1C", X"FD", --0640
  X"CB", X"01", X"7E", X"28", X"14", X"EF", X"F1", X"2B", --0648
  X"79", X"3D", X"B0", X"28", X"04", X"CD", X"AC", X"05", --0650
  X"24", X"1A", X"E6", X"DF", X"FE", X"50", X"C2", X"12", --0658
  X"19", X"2A", X"5D", X"5C", X"7E", X"FE", X"3B", X"C2", --0660
  X"12", X"19", X"EF", X"20", X"00", X"EF", X"82", X"1C", --0668
  X"FD", X"CB", X"01", X"7E", X"28", X"07", X"EF", X"99", --0670
  X"1E", X"ED", X"43", X"71", X"5B", X"EF", X"18", X"00", --0678
  X"FE", X"0D", X"28", X"05", X"FE", X"3A", X"C2", X"12", --0680
  X"19", X"CD", X"A1", X"18", X"ED", X"4B", X"71", X"5B", --0688
  X"78", X"B1", X"20", X"04", X"CD", X"AC", X"05", X"25", --0690
  X"21", X"B8", X"06", X"5E", X"23", X"56", X"23", X"EB", --0698
  X"7C", X"FE", X"25", X"30", X"0A", X"A7", X"ED", X"42", --06A0
  X"30", X"05", X"EB", X"23", X"23", X"18", X"EC", X"EB", --06A8
  X"5E", X"23", X"56", X"ED", X"53", X"5F", X"5B", X"C9", --06B0
  X"32", X"00", X"A5", X"0A", X"6E", X"00", X"D4", X"04", --06B8
  X"2C", X"01", X"C3", X"01", X"58", X"02", X"E0", X"00", --06C0
  X"B0", X"04", X"6E", X"00", X"60", X"09", X"36", X"00", --06C8
  X"C0", X"12", X"19", X"00", X"80", X"25", X"0B", X"00", --06D0
  X"21", X"61", X"5B", X"7E", X"A7", X"28", X"06", X"36", --06D8
  X"00", X"23", X"7E", X"37", X"C9", X"CD", X"D6", X"05", --06E0
  X"F3", X"D9", X"ED", X"5B", X"5F", X"5B", X"2A", X"5F", --06E8
  X"5B", X"CB", X"3C", X"CB", X"1D", X"B7", X"06", X"FA", --06F0
  X"D9", X"0E", X"FD", X"16", X"FF", X"1E", X"BF", X"42", --06F8
  X"3E", X"0E", X"ED", X"79", X"ED", X"78", X"F6", X"F0", --0700
  X"E6", X"FB", X"43", X"ED", X"79", X"67", X"42", X"ED", --0708
  X"78", X"E6", X"80", X"28", X"09", X"D9", X"05", X"D9", --0710
  X"20", X"F4", X"AF", X"F5", X"18", X"39", X"ED", X"78", --0718
  X"E6", X"80", X"20", X"F1", X"ED", X"78", X"E6", X"80", --0720
  X"20", X"EB", X"D9", X"01", X"FD", X"FF", X"3E", X"80", --0728
  X"08", X"19", X"00", X"00", X"00", X"00", X"2B", X"7C", --0730
  X"B5", X"20", X"FB", X"ED", X"78", X"E6", X"80", X"CA", --0738
  X"4B", X"07", X"08", X"37", X"1F", X"38", X"0D", X"08", --0740
  X"C3", X"31", X"07", X"08", X"B7", X"1F", X"38", X"04", --0748
  X"08", X"C3", X"31", X"07", X"37", X"F5", X"D9", X"7C", --0750
  X"F6", X"04", X"43", X"ED", X"79", X"D9", X"62", X"6B", --0758
  X"01", X"07", X"00", X"B7", X"ED", X"42", X"2B", X"7C", --0760
  X"B5", X"20", X"FB", X"01", X"FD", X"FF", X"19", X"19", --0768
  X"19", X"ED", X"78", X"E6", X"80", X"28", X"08", X"2B", --0770
  X"7C", X"B5", X"20", X"F5", X"F1", X"FB", X"C9", X"ED", --0778
  X"78", X"E6", X"80", X"20", X"EC", X"ED", X"78", X"E6", --0780
  X"80", X"20", X"E6", X"62", X"6B", X"01", X"02", X"00", --0788
  X"CB", X"3C", X"CB", X"1D", X"B7", X"ED", X"42", X"01", --0790
  X"FD", X"FF", X"3E", X"80", X"08", X"00", X"00", X"00", --0798
  X"00", X"19", X"2B", X"7C", X"B5", X"20", X"FB", X"ED", --07A0
  X"78", X"E6", X"80", X"CA", X"B7", X"07", X"08", X"37", --07A8
  X"1F", X"38", X"0D", X"08", X"C3", X"9D", X"07", X"08", --07B0
  X"B7", X"1F", X"38", X"04", X"08", X"C3", X"9D", X"07", --07B8
  X"21", X"61", X"5B", X"36", X"01", X"23", X"77", X"F1", --07C0
  X"FB", X"C9", X"F5", X"3A", X"65", X"5B", X"B7", X"28", --07C8
  X"0F", X"3D", X"32", X"65", X"5B", X"20", X"04", X"F1", --07D0
  X"C3", X"72", X"08", X"F1", X"32", X"0F", X"5C", X"C9", --07D8
  X"F1", X"FE", X"A3", X"38", X"0D", X"2A", X"5A", X"5B", --07E0
  X"E5", X"EF", X"52", X"0B", X"E1", X"22", X"5A", X"5B", --07E8
  X"37", X"C9", X"21", X"3B", X"5C", X"CB", X"86", X"FE", --07F0
  X"20", X"20", X"02", X"CB", X"C6", X"FE", X"7F", X"38", --07F8
  X"02", X"3E", X"3F", X"FE", X"20", X"38", X"17", X"F5", --0800
  X"21", X"63", X"5B", X"34", X"3A", X"64", X"5B", X"BE", --0808
  X"30", X"08", X"CD", X"22", X"08", X"3E", X"01", X"32", --0810
  X"63", X"5B", X"F1", X"C3", X"A3", X"08", X"FE", X"0D", --0818
  X"20", X"0E", X"AF", X"32", X"63", X"5B", X"3E", X"0D", --0820
  X"CD", X"A3", X"08", X"3E", X"0A", X"C3", X"A3", X"08", --0828
  X"FE", X"06", X"20", X"1F", X"ED", X"4B", X"63", X"5B", --0830
  X"1E", X"00", X"1C", X"0C", X"79", X"B8", X"28", X"08", --0838
  X"D6", X"08", X"28", X"04", X"30", X"FA", X"18", X"F2", --0840
  X"D5", X"3E", X"20", X"CD", X"CA", X"07", X"D1", X"1D", --0848
  X"C8", X"18", X"F5", X"FE", X"16", X"28", X"09", X"FE", --0850
  X"17", X"28", X"05", X"FE", X"10", X"D8", X"18", X"09", --0858
  X"32", X"0E", X"5C", X"3E", X"02", X"32", X"65", X"5B", --0860
  X"C9", X"32", X"0E", X"5C", X"3E", X"02", X"32", X"65", --0868
  X"5B", X"C9", X"57", X"3A", X"0E", X"5C", X"FE", X"16", --0870
  X"28", X"08", X"FE", X"17", X"3F", X"C0", X"3A", X"0F", --0878
  X"5C", X"57", X"3A", X"64", X"5B", X"BA", X"28", X"02", --0880
  X"30", X"06", X"47", X"7A", X"90", X"57", X"18", X"F2", --0888
  X"7A", X"B7", X"CA", X"22", X"08", X"3A", X"63", X"5B", --0890
  X"BA", X"C8", X"D5", X"3E", X"20", X"CD", X"CA", X"07", --0898
  X"D1", X"18", X"F2", X"F5", X"0E", X"FD", X"16", X"FF", --08A0
  X"1E", X"BF", X"42", X"3E", X"0E", X"ED", X"79", X"CD", --08A8
  X"D6", X"05", X"ED", X"78", X"E6", X"40", X"20", X"F7", --08B0
  X"2A", X"5F", X"5B", X"11", X"02", X"00", X"B7", X"ED", --08B8
  X"52", X"EB", X"F1", X"2F", X"37", X"06", X"0B", X"F3", --08C0
  X"C5", X"F5", X"3E", X"FE", X"62", X"6B", X"01", X"FD", --08C8
  X"BF", X"D2", X"DA", X"08", X"E6", X"F7", X"ED", X"79", --08D0
  X"18", X"06", X"F6", X"08", X"ED", X"79", X"18", X"00", --08D8
  X"2B", X"7C", X"B5", X"20", X"FB", X"00", X"00", X"00", --08E0
  X"F1", X"C1", X"B7", X"1F", X"10", X"DA", X"FB", X"C9", --08E8
  X"21", X"72", X"5B", X"36", X"2B", X"21", X"79", X"09", --08F0
  X"CD", X"5F", X"09", X"CD", X"15", X"09", X"21", X"80", --08F8
  X"09", X"CD", X"5F", X"09", X"21", X"72", X"5B", X"AF", --0900
  X"BE", X"28", X"03", X"35", X"18", X"E7", X"21", X"82", --0908
  X"09", X"CD", X"5F", X"09", X"C9", X"21", X"71", X"5B", --0910
  X"36", X"FF", X"CD", X"26", X"09", X"21", X"71", X"5B", --0918
  X"AF", X"BE", X"C8", X"35", X"18", X"F4", X"11", X"00", --0920
  X"C0", X"ED", X"4B", X"71", X"5B", X"37", X"CB", X"10", --0928
  X"37", X"CB", X"10", X"79", X"2F", X"4F", X"AF", X"F5", --0930
  X"D5", X"C5", X"CD", X"6D", X"09", X"C1", X"D1", X"1E", --0938
  X"00", X"28", X"01", X"5A", X"F1", X"B3", X"F5", X"05", --0940
  X"CB", X"3A", X"CB", X"3A", X"D5", X"C5", X"30", X"EA", --0948
  X"C1", X"D1", X"F1", X"06", X"03", X"C5", X"F5", X"CD", --0950
  X"A3", X"08", X"F1", X"C1", X"10", X"F7", X"C9", X"46", --0958
  X"23", X"7E", X"E5", X"C5", X"CD", X"A3", X"08", X"C1", --0960
  X"E1", X"23", X"10", X"F5", X"C9", X"EF", X"AA", X"22", --0968
  X"47", X"04", X"AF", X"37", X"1F", X"10", X"FD", X"A6", --0970
  X"C9", X"06", X"1B", X"31", X"1B", X"4C", X"00", X"03", --0978
  X"01", X"0A", X"02", X"1B", X"32", X"F3", X"C5", X"11", --0980
  X"37", X"00", X"21", X"3C", X"00", X"19", X"10", X"FD", --0988
  X"4D", X"44", X"EF", X"30", X"00", X"F3", X"D5", X"FD", --0990
  X"E1", X"E5", X"DD", X"E1", X"FD", X"36", X"10", X"FF", --0998
  X"01", X"C9", X"FF", X"DD", X"09", X"DD", X"36", X"03", --09A0
  X"3C", X"DD", X"36", X"01", X"FF", X"DD", X"36", X"04", --09A8
  X"0F", X"DD", X"36", X"05", X"05", X"DD", X"36", X"21", --09B0
  X"00", X"DD", X"36", X"0A", X"00", X"DD", X"36", X"0B", --09B8
  X"00", X"DD", X"36", X"16", X"FF", X"DD", X"36", X"17", --09C0
  X"00", X"DD", X"36", X"18", X"00", X"EF", X"F1", X"2B", --09C8
  X"F3", X"DD", X"73", X"06", X"DD", X"72", X"07", X"DD", --09D0
  X"73", X"0C", X"DD", X"72", X"0D", X"EB", X"09", X"DD", --09D8
  X"75", X"08", X"DD", X"74", X"09", X"C1", X"C5", X"05", --09E0
  X"48", X"06", X"00", X"CB", X"21", X"FD", X"E5", X"E1", --09E8
  X"09", X"DD", X"E5", X"C1", X"71", X"23", X"70", X"B7", --09F0
  X"FD", X"CB", X"10", X"16", X"C1", X"05", X"C5", X"DD", --09F8
  X"70", X"02", X"20", X"9C", X"C1", X"FD", X"36", X"27", --0A00
  X"1A", X"FD", X"36", X"28", X"0B", X"FD", X"E5", X"E1", --0A08
  X"01", X"2B", X"00", X"09", X"EB", X"21", X"31", X"0A", --0A10
  X"01", X"0D", X"00", X"ED", X"B0", X"16", X"07", X"1E", --0A18
  X"F8", X"CD", X"7C", X"0E", X"16", X"0B", X"1E", X"FF", --0A20
  X"CD", X"7C", X"0E", X"14", X"CD", X"7C", X"0E", X"18", --0A28
  X"4C", X"EF", X"A4", X"01", X"05", X"34", X"DF", X"75", --0A30
  X"F4", X"38", X"75", X"05", X"38", X"C9", X"3E", X"7F", --0A38
  X"DB", X"FE", X"1F", X"D8", X"3E", X"FE", X"DB", X"FE", --0A40
  X"1F", X"C9", X"01", X"11", X"00", X"18", X"03", X"01", --0A48
  X"00", X"00", X"FD", X"E5", X"E1", X"09", X"FD", X"75", --0A50
  X"23", X"FD", X"74", X"24", X"FD", X"7E", X"10", X"FD", --0A58
  X"77", X"22", X"FD", X"36", X"21", X"01", X"C9", X"5E", --0A60
  X"23", X"56", X"D5", X"DD", X"E1", X"C9", X"FD", X"6E", --0A68
  X"23", X"FD", X"66", X"24", X"23", X"23", X"FD", X"75", --0A70
  X"23", X"FD", X"74", X"24", X"C9", X"CD", X"4F", X"0A", --0A78
  X"FD", X"CB", X"22", X"1E", X"38", X"06", X"CD", X"67", --0A80
  X"0A", X"CD", X"5C", X"0B", X"FD", X"CB", X"21", X"26", --0A88
  X"38", X"05", X"CD", X"6E", X"0A", X"18", X"E9", X"CD", --0A90
  X"91", X"0F", X"D5", X"CD", X"42", X"0F", X"D1", X"FD", --0A98
  X"7E", X"10", X"FE", X"FF", X"20", X"05", X"CD", X"93", --0AA0
  X"0E", X"FB", X"C9", X"1B", X"CD", X"76", X"0F", X"CD", --0AA8
  X"C1", X"0F", X"CD", X"91", X"0F", X"18", X"E8", X"48", --0AB0
  X"5A", X"59", X"58", X"57", X"55", X"56", X"4D", X"54", --0AB8
  X"29", X"28", X"4E", X"4F", X"21", X"CD", X"E3", X"0E", --0AC0
  X"D8", X"DD", X"34", X"06", X"C0", X"DD", X"34", X"07", --0AC8
  X"C9", X"E5", X"0E", X"00", X"CD", X"C5", X"0A", X"38", --0AD0
  X"08", X"FE", X"26", X"20", X"0F", X"3E", X"80", X"E1", --0AD8
  X"C9", X"FD", X"7E", X"21", X"FD", X"B6", X"10", X"FD", --0AE0
  X"77", X"10", X"18", X"F3", X"FE", X"23", X"20", X"03", --0AE8
  X"0C", X"18", X"E1", X"FE", X"24", X"20", X"03", X"0D", --0AF0
  X"18", X"DA", X"CB", X"6F", X"20", X"06", X"F5", X"3E", --0AF8
  X"0C", X"81", X"4F", X"F1", X"E6", X"DF", X"D6", X"41", --0B00
  X"DA", X"22", X"0F", X"FE", X"07", X"D2", X"22", X"0F", --0B08
  X"C5", X"06", X"00", X"4F", X"21", X"F9", X"0D", X"09", --0B10
  X"7E", X"C1", X"81", X"E1", X"C9", X"E5", X"D5", X"DD", --0B18
  X"6E", X"06", X"DD", X"66", X"07", X"11", X"00", X"00", --0B20
  X"7E", X"FE", X"30", X"38", X"18", X"FE", X"3A", X"30", --0B28
  X"14", X"23", X"E5", X"CD", X"50", X"0B", X"D6", X"30", --0B30
  X"26", X"00", X"6F", X"19", X"38", X"04", X"EB", X"E1", --0B38
  X"18", X"E6", X"C3", X"1A", X"0F", X"DD", X"75", X"06", --0B40
  X"DD", X"74", X"07", X"D5", X"C1", X"D1", X"E1", X"C9", --0B48
  X"21", X"00", X"00", X"06", X"0A", X"19", X"38", X"EA", --0B50
  X"10", X"FB", X"EB", X"C9", X"CD", X"3E", X"0A", X"38", --0B58
  X"08", X"CD", X"93", X"0E", X"FB", X"CD", X"AC", X"05", --0B60
  X"14", X"CD", X"C5", X"0A", X"DA", X"A2", X"0D", X"CD", --0B68
  X"F0", X"0D", X"06", X"00", X"CB", X"21", X"21", X"CA", --0B70
  X"0D", X"09", X"5E", X"23", X"56", X"EB", X"CD", X"84", --0B78
  X"0B", X"18", X"D9", X"C9", X"E9", X"CD", X"C5", X"0A", --0B80
  X"DA", X"A1", X"0D", X"FE", X"21", X"C8", X"18", X"F5", --0B88
  X"CD", X"1D", X"0B", X"79", X"FE", X"09", X"D2", X"12", --0B90
  X"0F", X"CB", X"27", X"CB", X"27", X"47", X"CB", X"27", --0B98
  X"80", X"DD", X"77", X"03", X"C9", X"C9", X"DD", X"7E", --0BA0
  X"0B", X"3C", X"FE", X"05", X"CA", X"2A", X"0F", X"DD", --0BA8
  X"77", X"0B", X"11", X"0C", X"00", X"CD", X"27", X"0C", --0BB0
  X"DD", X"7E", X"06", X"77", X"23", X"DD", X"7E", X"07", --0BB8
  X"77", X"C9", X"DD", X"7E", X"16", X"11", X"17", X"00", --0BC0
  X"B7", X"FA", X"F0", X"0B", X"CD", X"27", X"0C", X"DD", --0BC8
  X"7E", X"06", X"BE", X"20", X"1B", X"23", X"DD", X"7E", --0BD0
  X"07", X"BE", X"20", X"14", X"DD", X"35", X"16", X"DD", --0BD8
  X"7E", X"16", X"B7", X"F0", X"DD", X"CB", X"0A", X"46", --0BE0
  X"C8", X"DD", X"36", X"16", X"00", X"AF", X"18", X"1B", --0BE8
  X"DD", X"7E", X"16", X"3C", X"FE", X"05", X"CA", X"2A", --0BF0
  X"0F", X"DD", X"77", X"16", X"CD", X"27", X"0C", X"DD", --0BF8
  X"7E", X"06", X"77", X"23", X"DD", X"7E", X"07", X"77", --0C00
  X"DD", X"7E", X"0B", X"11", X"0C", X"00", X"CD", X"27", --0C08
  X"0C", X"7E", X"DD", X"77", X"06", X"23", X"7E", X"DD", --0C10
  X"77", X"07", X"DD", X"35", X"0B", X"F0", X"DD", X"36", --0C18
  X"0B", X"00", X"DD", X"CB", X"0A", X"C6", X"C9", X"DD", --0C20
  X"E5", X"E1", X"19", X"06", X"00", X"4F", X"CB", X"21", --0C28
  X"09", X"C9", X"CD", X"1D", X"0B", X"78", X"B7", X"C2", --0C30
  X"12", X"0F", X"79", X"FE", X"3C", X"DA", X"12", X"0F", --0C38
  X"FE", X"F1", X"D2", X"12", X"0F", X"DD", X"7E", X"02", --0C40
  X"B7", X"C0", X"06", X"00", X"C5", X"E1", X"29", X"29", --0C48
  X"E5", X"C1", X"FD", X"E5", X"EF", X"2B", X"2D", X"F3", --0C50
  X"FD", X"E1", X"FD", X"E5", X"FD", X"E5", X"E1", X"01", --0C58
  X"2B", X"00", X"09", X"FD", X"21", X"3A", X"5C", X"E5", --0C60
  X"21", X"76", X"0C", X"22", X"5A", X"5B", X"21", X"14", --0C68
  X"5B", X"E3", X"E5", X"C3", X"00", X"5B", X"F3", X"EF", --0C70
  X"A2", X"2D", X"F3", X"FD", X"E1", X"FD", X"71", X"27", --0C78
  X"FD", X"70", X"28", X"C9", X"CD", X"1D", X"0B", X"79", --0C80
  X"FE", X"40", X"D2", X"12", X"0F", X"2F", X"5F", X"16", --0C88
  X"07", X"CD", X"7C", X"0E", X"C9", X"CD", X"1D", X"0B", --0C90
  X"79", X"FE", X"10", X"D2", X"12", X"0F", X"DD", X"77", --0C98
  X"04", X"DD", X"5E", X"02", X"3E", X"08", X"83", X"57", --0CA0
  X"59", X"CD", X"7C", X"0E", X"C9", X"DD", X"5E", X"02", --0CA8
  X"3E", X"08", X"83", X"57", X"1E", X"1F", X"DD", X"73", --0CB0
  X"04", X"C9", X"CD", X"1D", X"0B", X"79", X"FE", X"08", --0CB8
  X"D2", X"12", X"0F", X"06", X"00", X"21", X"E8", X"0D", --0CC0
  X"09", X"7E", X"FD", X"77", X"29", X"C9", X"CD", X"1D", --0CC8
  X"0B", X"16", X"0B", X"59", X"CD", X"7C", X"0E", X"14", --0CD0
  X"58", X"CD", X"7C", X"0E", X"C9", X"CD", X"1D", X"0B", --0CD8
  X"79", X"3D", X"FA", X"12", X"0F", X"FE", X"10", X"D2", --0CE0
  X"12", X"0F", X"DD", X"77", X"01", X"C9", X"CD", X"1D", --0CE8
  X"0B", X"79", X"CD", X"A3", X"11", X"C9", X"FD", X"36", --0CF0
  X"10", X"FF", X"C9", X"CD", X"19", X"0E", X"DA", X"81", --0CF8
  X"0D", X"CD", X"AC", X"0D", X"CD", X"B4", X"0D", X"AF", --0D00
  X"DD", X"77", X"21", X"CD", X"C8", X"0E", X"CD", X"1D", --0D08
  X"0B", X"79", X"B7", X"CA", X"12", X"0F", X"FE", X"0D", --0D10
  X"D2", X"12", X"0F", X"FE", X"0A", X"38", X"13", X"CD", --0D18
  X"00", X"0E", X"CD", X"74", X"0D", X"73", X"23", X"72", --0D20
  X"CD", X"74", X"0D", X"23", X"73", X"23", X"72", X"23", --0D28
  X"18", X"06", X"DD", X"71", X"05", X"CD", X"00", X"0E", --0D30
  X"CD", X"74", X"0D", X"CD", X"E3", X"0E", X"FE", X"5F", --0D38
  X"20", X"2C", X"CD", X"C5", X"0A", X"CD", X"1D", X"0B", --0D40
  X"79", X"FE", X"0A", X"38", X"12", X"E5", X"D5", X"CD", --0D48
  X"00", X"0E", X"E1", X"19", X"4B", X"42", X"EB", X"E1", --0D50
  X"73", X"23", X"72", X"59", X"50", X"18", X"C9", X"DD", --0D58
  X"71", X"05", X"E5", X"D5", X"CD", X"00", X"0E", X"E1", --0D60
  X"19", X"EB", X"E1", X"C3", X"3B", X"0D", X"73", X"23", --0D68
  X"72", X"C3", X"9C", X"0D", X"DD", X"7E", X"21", X"3C", --0D70
  X"FE", X"0B", X"CA", X"3A", X"0F", X"DD", X"77", X"21", --0D78
  X"C9", X"CD", X"C8", X"0E", X"DD", X"36", X"21", X"01", --0D80
  X"CD", X"AC", X"0D", X"CD", X"B4", X"0D", X"DD", X"4E", --0D88
  X"05", X"E5", X"CD", X"00", X"0E", X"E1", X"73", X"23", --0D90
  X"72", X"C3", X"9C", X"0D", X"E1", X"23", X"23", X"E5", --0D98
  X"C9", X"E1", X"FD", X"7E", X"21", X"FD", X"B6", X"10", --0DA0
  X"FD", X"77", X"10", X"C9", X"DD", X"E5", X"E1", X"01", --0DA8
  X"22", X"00", X"09", X"C9", X"E5", X"FD", X"E5", X"E1", --0DB0
  X"01", X"11", X"00", X"09", X"06", X"00", X"DD", X"4E", --0DB8
  X"02", X"CB", X"21", X"09", X"D1", X"73", X"23", X"72", --0DC0
  X"EB", X"C9", X"FB", X"0C", X"85", X"0B", X"90", X"0B", --0DC8
  X"A5", X"0B", X"A6", X"0B", X"C2", X"0B", X"32", X"0C", --0DD0
  X"84", X"0C", X"95", X"0C", X"AD", X"0C", X"BA", X"0C", --0DD8
  X"CE", X"0C", X"DD", X"0C", X"EE", X"0C", X"F6", X"0C", --0DE0
  X"00", X"04", X"0B", X"0D", X"08", X"0C", X"0E", X"0A", --0DE8
  X"01", X"0F", X"00", X"21", X"B7", X"0A", X"ED", X"B1", --0DF0
  X"C9", X"09", X"0B", X"00", X"02", X"04", X"05", X"07", --0DF8
  X"E5", X"06", X"00", X"21", X"0C", X"0E", X"09", X"16", --0E00
  X"00", X"5E", X"E1", X"C9", X"80", X"06", X"09", X"0C", --0E08
  X"12", X"18", X"24", X"30", X"48", X"60", X"04", X"08", --0E10
  X"10", X"FE", X"30", X"D8", X"FE", X"3A", X"3F", X"C9", --0E18
  X"4F", X"DD", X"7E", X"03", X"81", X"FE", X"80", X"D2", --0E20
  X"32", X"0F", X"4F", X"DD", X"7E", X"02", X"B7", X"20", --0E28
  X"0E", X"79", X"2F", X"E6", X"7F", X"CB", X"3F", X"CB", --0E30
  X"3F", X"16", X"06", X"5F", X"CD", X"7C", X"0E", X"DD", --0E38
  X"71", X"00", X"DD", X"7E", X"02", X"FE", X"03", X"D0", --0E40
  X"21", X"96", X"10", X"06", X"00", X"79", X"D6", X"15", --0E48
  X"30", X"05", X"11", X"BF", X"0F", X"18", X"07", X"4F", --0E50
  X"CB", X"21", X"09", X"5E", X"23", X"56", X"EB", X"DD", --0E58
  X"56", X"02", X"CB", X"22", X"5D", X"CD", X"7C", X"0E", --0E60
  X"14", X"5C", X"CD", X"7C", X"0E", X"DD", X"CB", X"04", --0E68
  X"66", X"C8", X"16", X"0D", X"FD", X"7E", X"29", X"5F", --0E70
  X"CD", X"7C", X"0E", X"C9", X"C5", X"01", X"FD", X"FF", --0E78
  X"ED", X"51", X"01", X"FD", X"BF", X"ED", X"59", X"C1", --0E80
  X"C9", X"C5", X"01", X"FD", X"FF", X"ED", X"79", X"ED", --0E88
  X"78", X"C1", X"C9", X"16", X"07", X"1E", X"FF", X"CD", --0E90
  X"7C", X"0E", X"16", X"08", X"1E", X"00", X"CD", X"7C", --0E98
  X"0E", X"14", X"CD", X"7C", X"0E", X"14", X"CD", X"7C", --0EA0
  X"0E", X"CD", X"4F", X"0A", X"FD", X"CB", X"22", X"1E", --0EA8
  X"38", X"06", X"CD", X"67", X"0A", X"CD", X"8D", X"11", --0EB0
  X"FD", X"CB", X"21", X"26", X"38", X"05", X"CD", X"6E", --0EB8
  X"0A", X"18", X"E9", X"FD", X"21", X"3A", X"5C", X"C9", --0EC0
  X"E5", X"D5", X"DD", X"6E", X"06", X"DD", X"66", X"07", --0EC8
  X"2B", X"7E", X"FE", X"20", X"28", X"FA", X"FE", X"0D", --0ED0
  X"28", X"F6", X"DD", X"75", X"06", X"DD", X"74", X"07", --0ED8
  X"D1", X"E1", X"C9", X"E5", X"D5", X"C5", X"DD", X"6E", --0EE0
  X"06", X"DD", X"66", X"07", X"7C", X"DD", X"BE", X"09", --0EE8
  X"20", X"09", X"7D", X"DD", X"BE", X"08", X"20", X"03", --0EF0
  X"37", X"18", X"0A", X"7E", X"FE", X"20", X"28", X"09", --0EF8
  X"FE", X"0D", X"28", X"05", X"B7", X"C1", X"D1", X"E1", --0F00
  X"C9", X"23", X"DD", X"75", X"06", X"DD", X"74", X"07", --0F08
  X"18", X"DA", X"CD", X"93", X"0E", X"FB", X"CD", X"AC", --0F10
  X"05", X"29", X"CD", X"93", X"0E", X"FB", X"CD", X"AC", --0F18
  X"05", X"27", X"CD", X"93", X"0E", X"FB", X"CD", X"AC", --0F20
  X"05", X"26", X"CD", X"93", X"0E", X"FB", X"CD", X"AC", --0F28
  X"05", X"1F", X"CD", X"93", X"0E", X"FB", X"CD", X"AC", --0F30
  X"05", X"28", X"CD", X"93", X"0E", X"FB", X"CD", X"AC", --0F38
  X"05", X"2A", X"CD", X"4F", X"0A", X"FD", X"CB", X"22", --0F40
  X"1E", X"38", X"21", X"CD", X"67", X"0A", X"CD", X"D1", --0F48
  X"0A", X"FE", X"80", X"28", X"17", X"CD", X"20", X"0E", --0F50
  X"DD", X"7E", X"02", X"FE", X"03", X"30", X"0A", X"16", --0F58
  X"08", X"82", X"57", X"DD", X"5E", X"04", X"CD", X"7C", --0F60
  X"0E", X"CD", X"6E", X"11", X"FD", X"CB", X"21", X"26", --0F68
  X"D8", X"CD", X"6E", X"0A", X"18", X"CF", X"E5", X"FD", --0F70
  X"6E", X"27", X"FD", X"66", X"28", X"01", X"64", X"00", --0F78
  X"B7", X"ED", X"42", X"E5", X"C1", X"E1", X"0B", X"78", --0F80
  X"B1", X"20", X"FB", X"1B", X"7A", X"B3", X"20", X"E6", --0F88
  X"C9", X"11", X"FF", X"FF", X"CD", X"4A", X"0A", X"FD", --0F90
  X"CB", X"22", X"1E", X"38", X"12", X"D5", X"5E", X"23", --0F98
  X"56", X"EB", X"5E", X"23", X"56", X"D5", X"E1", X"C1", --0FA0
  X"B7", X"ED", X"42", X"38", X"02", X"C5", X"D1", X"FD", --0FA8
  X"CB", X"21", X"26", X"38", X"05", X"CD", X"6E", X"0A", --0FB0
  X"18", X"DD", X"FD", X"73", X"25", X"FD", X"72", X"26", --0FB8
  X"C9", X"AF", X"FD", X"77", X"2A", X"CD", X"4F", X"0A", --0FC0
  X"FD", X"CB", X"22", X"1E", X"DA", X"5A", X"10", X"CD", --0FC8
  X"67", X"0A", X"FD", X"E5", X"E1", X"01", X"11", X"00", --0FD0
  X"09", X"06", X"00", X"DD", X"4E", X"02", X"CB", X"21", --0FD8
  X"09", X"5E", X"23", X"56", X"EB", X"E5", X"5E", X"23", --0FE0
  X"56", X"EB", X"FD", X"5E", X"25", X"FD", X"56", X"26", --0FE8
  X"B7", X"ED", X"52", X"EB", X"E1", X"28", X"05", X"73", --0FF0
  X"23", X"72", X"18", X"5E", X"DD", X"7E", X"02", X"FE", --0FF8
  X"03", X"30", X"09", X"16", X"08", X"82", X"57", X"1E", --1000
  X"00", X"CD", X"7C", X"0E", X"CD", X"8D", X"11", X"DD", --1008
  X"E5", X"E1", X"01", X"21", X"00", X"09", X"35", X"20", --1010
  X"0D", X"CD", X"5C", X"0B", X"FD", X"7E", X"21", X"FD", --1018
  X"A6", X"10", X"20", X"36", X"18", X"17", X"FD", X"E5", --1020
  X"E1", X"01", X"11", X"00", X"09", X"06", X"00", X"DD", --1028
  X"4E", X"02", X"CB", X"21", X"09", X"5E", X"23", X"56", --1030
  X"13", X"13", X"72", X"2B", X"73", X"CD", X"D1", X"0A", --1038
  X"4F", X"FD", X"7E", X"21", X"FD", X"A6", X"10", X"20", --1040
  X"11", X"79", X"FE", X"80", X"28", X"0C", X"CD", X"20", --1048
  X"0E", X"FD", X"7E", X"21", X"FD", X"B6", X"2A", X"FD", --1050
  X"77", X"2A", X"FD", X"CB", X"21", X"26", X"38", X"06", --1058
  X"CD", X"6E", X"0A", X"C3", X"C8", X"0F", X"11", X"01", --1060
  X"00", X"CD", X"76", X"0F", X"CD", X"4F", X"0A", X"FD", --1068
  X"CB", X"2A", X"1E", X"30", X"17", X"CD", X"67", X"0A", --1070
  X"DD", X"7E", X"02", X"FE", X"03", X"30", X"0A", X"16", --1078
  X"08", X"82", X"57", X"DD", X"5E", X"04", X"CD", X"7C", --1080
  X"0E", X"CD", X"6E", X"11", X"FD", X"CB", X"21", X"26", --1088
  X"D8", X"CD", X"6E", X"0A", X"18", X"D9", X"BF", X"0F", --1090
  X"DC", X"0E", X"07", X"0E", X"3D", X"0D", X"7F", X"0C", --1098
  X"CC", X"0B", X"22", X"0B", X"82", X"0A", X"EB", X"09", --10A0
  X"5D", X"09", X"D6", X"08", X"57", X"08", X"DF", X"07", --10A8
  X"6E", X"07", X"03", X"07", X"9F", X"06", X"40", X"06", --10B0
  X"E6", X"05", X"91", X"05", X"41", X"05", X"F6", X"04", --10B8
  X"AE", X"04", X"6B", X"04", X"2C", X"04", X"F0", X"03", --10C0
  X"B7", X"03", X"82", X"03", X"4F", X"03", X"20", X"03", --10C8
  X"F3", X"02", X"C8", X"02", X"A1", X"02", X"7B", X"02", --10D0
  X"57", X"02", X"36", X"02", X"16", X"02", X"F8", X"01", --10D8
  X"DC", X"01", X"C1", X"01", X"A8", X"01", X"90", X"01", --10E0
  X"79", X"01", X"64", X"01", X"50", X"01", X"3D", X"01", --10E8
  X"2C", X"01", X"1B", X"01", X"0B", X"01", X"FC", X"00", --10F0
  X"EE", X"00", X"E0", X"00", X"D4", X"00", X"C8", X"00", --10F8
  X"BD", X"00", X"B2", X"00", X"A8", X"00", X"9F", X"00", --1100
  X"96", X"00", X"8D", X"00", X"85", X"00", X"7E", X"00", --1108
  X"77", X"00", X"70", X"00", X"6A", X"00", X"64", X"00", --1110
  X"5E", X"00", X"59", X"00", X"54", X"00", X"4F", X"00", --1118
  X"4B", X"00", X"47", X"00", X"43", X"00", X"3F", X"00", --1120
  X"3B", X"00", X"38", X"00", X"35", X"00", X"32", X"00", --1128
  X"2F", X"00", X"2D", X"00", X"2A", X"00", X"28", X"00", --1130
  X"25", X"00", X"23", X"00", X"21", X"00", X"1F", X"00", --1138
  X"1E", X"00", X"1C", X"00", X"1A", X"00", X"19", X"00", --1140
  X"18", X"00", X"16", X"00", X"15", X"00", X"14", X"00", --1148
  X"13", X"00", X"12", X"00", X"11", X"00", X"10", X"00", --1150
  X"0F", X"00", X"0E", X"00", X"0D", X"00", X"0C", X"00", --1158
  X"0C", X"00", X"0B", X"00", X"0B", X"00", X"0A", X"00", --1160
  X"09", X"00", X"09", X"00", X"08", X"00", X"DD", X"7E", --1168
  X"01", X"B7", X"F8", X"F6", X"90", X"CD", X"A3", X"11", --1170
  X"DD", X"7E", X"00", X"CD", X"A3", X"11", X"DD", X"7E", --1178
  X"04", X"CB", X"A7", X"CB", X"27", X"CB", X"27", X"CB", --1180
  X"27", X"CD", X"A3", X"11", X"C9", X"DD", X"7E", X"01", --1188
  X"B7", X"F8", X"F6", X"80", X"CD", X"A3", X"11", X"DD", --1190
  X"7E", X"00", X"CD", X"A3", X"11", X"3E", X"40", X"CD", --1198
  X"A3", X"11", X"C9", X"6F", X"01", X"FD", X"FF", X"3E", --11A0
  X"0E", X"ED", X"79", X"01", X"FD", X"BF", X"3E", X"FA", --11A8
  X"ED", X"79", X"1E", X"03", X"1D", X"20", X"FD", X"00", --11B0
  X"00", X"00", X"00", X"7D", X"16", X"08", X"1F", X"6F", --11B8
  X"D2", X"C9", X"11", X"3E", X"FE", X"ED", X"79", X"18", --11C0
  X"06", X"3E", X"FA", X"ED", X"79", X"18", X"00", X"1E", --11C8
  X"02", X"1D", X"20", X"FD", X"00", X"C6", X"00", X"7D", --11D0
  X"15", X"20", X"E3", X"00", X"00", X"C6", X"00", X"00", --11D8
  X"00", X"3E", X"FE", X"ED", X"79", X"1E", X"06", X"1D", --11E0
  X"20", X"FD", X"C9", X"21", X"66", X"5B", X"CB", X"EE", --11E8
  X"18", X"13", X"21", X"66", X"5B", X"CB", X"E6", X"18", --11F0
  X"0C", X"21", X"66", X"5B", X"CB", X"FE", X"18", X"05", --11F8
  X"21", X"66", X"5B", X"CB", X"F6", X"21", X"66", X"5B", --1200
  X"CB", X"9E", X"DF", X"FE", X"21", X"C2", X"BE", X"13", --1208
  X"21", X"66", X"5B", X"CB", X"DE", X"E7", X"C3", X"BE", --1210
  X"13", X"CD", X"AC", X"05", X"0B", X"22", X"74", X"5B", --1218
  X"DD", X"7E", X"00", X"32", X"71", X"5B", X"DD", X"6E", --1220
  X"0B", X"DD", X"66", X"0C", X"22", X"72", X"5B", X"DD", --1228
  X"6E", X"0D", X"DD", X"66", X"0E", X"22", X"78", X"5B", --1230
  X"DD", X"6E", X"0F", X"DD", X"66", X"10", X"22", X"76", --1238
  X"5B", X"B7", X"28", X"0A", X"FE", X"03", X"28", X"06", --1240
  X"DD", X"7E", X"0E", X"32", X"76", X"5B", X"DD", X"E5", --1248
  X"E1", X"23", X"11", X"67", X"5B", X"01", X"0A", X"00", --1250
  X"ED", X"B0", X"21", X"66", X"5B", X"CB", X"6E", X"C2", --1258
  X"AD", X"1B", X"21", X"71", X"5B", X"11", X"7A", X"5B", --1260
  X"01", X"07", X"00", X"ED", X"B0", X"CD", X"2E", X"1C", --1268
  X"3A", X"7A", X"5B", X"47", X"3A", X"71", X"5B", X"B8", --1270
  X"20", X"06", X"FE", X"03", X"28", X"12", X"38", X"04", --1278
  X"CD", X"AC", X"05", X"1D", X"3A", X"66", X"5B", X"CB", --1280
  X"77", X"20", X"3A", X"CB", X"7F", X"CA", X"DB", X"12", --1288
  X"3A", X"66", X"5B", X"CB", X"77", X"28", X"04", X"CD", --1290
  X"AC", X"05", X"1C", X"2A", X"7B", X"5B", X"ED", X"5B", --1298
  X"72", X"5B", X"7C", X"B5", X"28", X"08", X"ED", X"52", --12A0
  X"30", X"04", X"CD", X"AC", X"05", X"1E", X"2A", X"7D", --12A8
  X"5B", X"7C", X"B5", X"20", X"03", X"2A", X"74", X"5B", --12B0
  X"3A", X"71", X"5B", X"A7", X"20", X"03", X"2A", X"53", --12B8
  X"5C", X"CD", X"7E", X"13", X"C9", X"ED", X"4B", X"72", --12C0
  X"5B", X"C5", X"03", X"EF", X"30", X"00", X"36", X"80", --12C8
  X"EB", X"D1", X"E5", X"CD", X"7E", X"13", X"E1", X"EF", --12D0
  X"CE", X"08", X"C9", X"ED", X"5B", X"72", X"5B", X"2A", --12D8
  X"7D", X"5B", X"E5", X"7C", X"B5", X"20", X"06", X"13", --12E0
  X"13", X"13", X"EB", X"18", X"09", X"2A", X"7B", X"5B", --12E8
  X"EB", X"37", X"ED", X"52", X"38", X"09", X"11", X"05", --12F0
  X"00", X"19", X"44", X"4D", X"EF", X"05", X"1F", X"E1", --12F8
  X"3A", X"71", X"5B", X"A7", X"28", X"2F", X"7C", X"B5", --1300
  X"28", X"0B", X"2B", X"46", X"2B", X"4E", X"2B", X"03", --1308
  X"03", X"03", X"EF", X"E8", X"19", X"2A", X"59", X"5C", --1310
  X"2B", X"ED", X"4B", X"72", X"5B", X"C5", X"03", X"03", --1318
  X"03", X"3A", X"7F", X"5B", X"F5", X"EF", X"55", X"16", --1320
  X"23", X"F1", X"77", X"D1", X"23", X"73", X"23", X"72", --1328
  X"23", X"CD", X"7E", X"13", X"C9", X"21", X"66", X"5B", --1330
  X"CB", X"8E", X"ED", X"5B", X"53", X"5C", X"2A", X"59", --1338
  X"5C", X"2B", X"EF", X"E5", X"19", X"ED", X"4B", X"72", --1340
  X"5B", X"2A", X"53", X"5C", X"EF", X"55", X"16", X"23", --1348
  X"ED", X"4B", X"76", X"5B", X"09", X"22", X"4B", X"5C", --1350
  X"3A", X"79", X"5B", X"67", X"E6", X"C0", X"20", X"10", --1358
  X"3A", X"78", X"5B", X"6F", X"22", X"42", X"5C", X"FD", --1360
  X"36", X"0A", X"00", X"21", X"66", X"5B", X"CB", X"CE", --1368
  X"2A", X"53", X"5C", X"ED", X"5B", X"72", X"5B", X"2B", --1370
  X"22", X"57", X"5C", X"23", X"18", X"B3", X"7A", X"B3", --1378
  X"C8", X"CD", X"4B", X"1C", X"C9", X"EF", X"8C", X"1C", --1380
  X"FD", X"CB", X"01", X"7E", X"C8", X"F5", X"EF", X"F1", --1388
  X"2B", X"F1", X"C9", X"E7", X"CD", X"85", X"13", X"C8", --1390
  X"F5", X"79", X"B0", X"28", X"1D", X"21", X"0A", X"00", --1398
  X"ED", X"42", X"38", X"16", X"D5", X"C5", X"21", X"67", --13A0
  X"5B", X"06", X"0A", X"3E", X"20", X"77", X"23", X"10", --13A8
  X"FC", X"C1", X"E1", X"11", X"67", X"5B", X"ED", X"B0", --13B0
  X"F1", X"C9", X"CD", X"AC", X"05", X"21", X"EF", X"8C", --13B8
  X"1C", X"FD", X"CB", X"01", X"7E", X"28", X"40", X"01", --13C0
  X"11", X"00", X"3A", X"74", X"5C", X"A7", X"28", X"02", --13C8
  X"0E", X"22", X"EF", X"30", X"00", X"D5", X"DD", X"E1", --13D0
  X"06", X"0B", X"3E", X"20", X"12", X"13", X"10", X"FC", --13D8
  X"DD", X"36", X"01", X"FF", X"EF", X"F1", X"2B", X"21", --13E0
  X"F6", X"FF", X"0B", X"09", X"03", X"30", X"11", X"3A", --13E8
  X"74", X"5C", X"A7", X"20", X"04", X"CD", X"AC", X"05", --13F0
  X"0E", X"78", X"B1", X"28", X"0A", X"01", X"0A", X"00", --13F8
  X"DD", X"E5", X"E1", X"23", X"EB", X"ED", X"B0", X"DF", --1400
  X"FE", X"E4", X"20", X"53", X"3A", X"74", X"5C", X"FE", --1408
  X"03", X"CA", X"19", X"12", X"E7", X"EF", X"B2", X"28", --1410
  X"30", X"15", X"21", X"00", X"00", X"FD", X"CB", X"01", --1418
  X"76", X"28", X"02", X"CB", X"F9", X"3A", X"74", X"5C", --1420
  X"3D", X"28", X"19", X"CD", X"AC", X"05", X"01", X"C2", --1428
  X"19", X"12", X"FD", X"CB", X"01", X"7E", X"28", X"19", --1430
  X"4E", X"23", X"7E", X"DD", X"77", X"0B", X"23", X"7E", --1438
  X"DD", X"77", X"0C", X"23", X"DD", X"71", X"0E", X"3E", --1440
  X"01", X"CB", X"71", X"28", X"01", X"3C", X"DD", X"77", --1448
  X"00", X"EB", X"E7", X"FE", X"29", X"20", X"D8", X"E7", --1450
  X"CD", X"A1", X"18", X"EB", X"C3", X"19", X"15", X"FE", --1458
  X"AA", X"20", X"1F", X"3A", X"74", X"5C", X"FE", X"03", --1460
  X"CA", X"19", X"12", X"E7", X"CD", X"A1", X"18", X"DD", --1468
  X"36", X"0B", X"00", X"DD", X"36", X"0C", X"1B", X"21", --1470
  X"00", X"40", X"DD", X"75", X"0D", X"DD", X"74", X"0E", --1478
  X"18", X"4D", X"FE", X"AF", X"20", X"4F", X"3A", X"74", --1480
  X"5C", X"FE", X"03", X"CA", X"19", X"12", X"E7", X"EF", --1488
  X"48", X"20", X"20", X"0C", X"3A", X"74", X"5C", X"A7", --1490
  X"CA", X"19", X"12", X"EF", X"E6", X"1C", X"18", X"0F", --1498
  X"EF", X"82", X"1C", X"DF", X"FE", X"2C", X"28", X"0C", --14A0
  X"3A", X"74", X"5C", X"A7", X"CA", X"19", X"12", X"EF", --14A8
  X"E6", X"1C", X"18", X"04", X"E7", X"EF", X"82", X"1C", --14B0
  X"CD", X"A1", X"18", X"EF", X"99", X"1E", X"DD", X"71", --14B8
  X"0B", X"DD", X"70", X"0C", X"EF", X"99", X"1E", X"DD", --14C0
  X"71", X"0D", X"DD", X"70", X"0E", X"60", X"69", X"DD", --14C8
  X"36", X"00", X"03", X"18", X"44", X"FE", X"CA", X"28", --14D0
  X"09", X"CD", X"A1", X"18", X"DD", X"36", X"0E", X"80", --14D8
  X"18", X"17", X"3A", X"74", X"5C", X"A7", X"C2", X"19", --14E0
  X"12", X"E7", X"EF", X"82", X"1C", X"CD", X"A1", X"18", --14E8
  X"EF", X"99", X"1E", X"DD", X"71", X"0D", X"DD", X"70", --14F0
  X"0E", X"DD", X"36", X"00", X"00", X"2A", X"59", X"5C", --14F8
  X"ED", X"5B", X"53", X"5C", X"37", X"ED", X"52", X"DD", --1500
  X"75", X"0B", X"DD", X"74", X"0C", X"2A", X"4B", X"5C", --1508
  X"ED", X"52", X"DD", X"75", X"0F", X"DD", X"74", X"10", --1510
  X"EB", X"3A", X"66", X"5B", X"CB", X"5F", X"C2", X"1D", --1518
  X"12", X"3A", X"74", X"5C", X"A7", X"20", X"04", X"EF", --1520
  X"70", X"09", X"C9", X"EF", X"61", X"07", X"C9", X"21", --1528
  X"F5", X"EE", X"CB", X"86", X"CB", X"CE", X"2A", X"49", --1530
  X"5C", X"7C", X"B5", X"20", X"03", X"22", X"06", X"EC", --1538
  X"3A", X"DB", X"F9", X"F5", X"2A", X"9A", X"FC", X"CD", --1540
  X"4A", X"33", X"22", X"D7", X"F9", X"CD", X"22", X"32", --1548
  X"CD", X"D6", X"30", X"F1", X"B7", X"28", X"0C", X"F5", --1550
  X"CD", X"DF", X"30", X"EB", X"CD", X"6A", X"32", X"F1", --1558
  X"3D", X"18", X"F1", X"0E", X"00", X"CD", X"B4", X"30", --1560
  X"41", X"3A", X"15", X"EC", X"4F", X"C5", X"D5", X"CD", --1568
  X"DF", X"30", X"3A", X"F5", X"EE", X"CB", X"4F", X"28", --1570
  X"1D", X"D5", X"E5", X"11", X"20", X"00", X"19", X"CB", --1578
  X"46", X"28", X"11", X"23", X"56", X"23", X"5E", X"B7", --1580
  X"2A", X"49", X"5C", X"ED", X"52", X"20", X"05", X"21", --1588
  X"F5", X"EE", X"CB", X"C6", X"E1", X"D1", X"C5", X"E5", --1590
  X"01", X"23", X"00", X"ED", X"B0", X"E1", X"C1", X"D5", --1598
  X"C5", X"EB", X"21", X"F5", X"EE", X"CB", X"46", X"28", --15A0
  X"2A", X"06", X"00", X"2A", X"06", X"EC", X"7C", X"B5", --15A8
  X"28", X"0E", X"E5", X"CD", X"41", X"2E", X"E1", X"30", --15B0
  X"12", X"2B", X"04", X"22", X"06", X"EC", X"18", X"EB", --15B8
  X"CD", X"41", X"2E", X"D4", X"63", X"2E", X"21", X"F5", --15C0
  X"EE", X"36", X"00", X"78", X"C1", X"C5", X"48", X"47", --15C8
  X"CD", X"11", X"2A", X"C1", X"D1", X"79", X"04", X"B8", --15D0
  X"30", X"95", X"3A", X"F5", X"EE", X"CB", X"4F", X"28", --15D8
  X"21", X"CB", X"47", X"20", X"1D", X"2A", X"49", X"5C", --15E0
  X"7C", X"B5", X"28", X"08", X"22", X"9A", X"FC", X"CD", --15E8
  X"22", X"32", X"18", X"09", X"22", X"9A", X"FC", X"CD", --15F0
  X"52", X"33", X"22", X"49", X"5C", X"D1", X"C1", X"C3", --15F8
  X"36", X"15", X"D1", X"C1", X"BF", X"F5", X"79", X"48", --1600
  X"CD", X"B4", X"30", X"EB", X"F5", X"CD", X"04", X"36", --1608
  X"F1", X"11", X"23", X"00", X"19", X"0C", X"B9", X"30", --1610
  X"F3", X"F1", X"C8", X"CD", X"07", X"2A", X"CD", X"78", --1618
  X"2B", X"2A", X"06", X"EC", X"2B", X"7C", X"B5", X"22", --1620
  X"06", X"EC", X"20", X"F2", X"C3", X"11", X"2A", X"C9", --1628
  X"06", X"00", X"3A", X"15", X"EC", X"57", X"C3", X"5E", --1630
  X"3B", X"06", X"00", X"E5", X"48", X"CD", X"B4", X"30", --1638
  X"CD", X"6A", X"32", X"E1", X"D0", X"CD", X"DF", X"30", --1640
  X"C5", X"E5", X"21", X"23", X"00", X"19", X"3A", X"15", --1648
  X"EC", X"4F", X"B8", X"28", X"0E", X"C5", X"C5", X"01", --1650
  X"23", X"00", X"ED", X"B0", X"C1", X"79", X"04", X"B8", --1658
  X"20", X"F4", X"C1", X"E1", X"CD", X"18", X"36", X"01", --1660
  X"23", X"00", X"ED", X"B0", X"37", X"C1", X"C9", X"06", --1668
  X"00", X"CD", X"2B", X"32", X"D0", X"C5", X"E5", X"3A", --1670
  X"15", X"EC", X"4F", X"CD", X"B4", X"30", X"CD", X"1E", --1678
  X"31", X"30", X"26", X"1B", X"21", X"23", X"00", X"19", --1680
  X"EB", X"C5", X"78", X"B9", X"28", X"0C", X"C5", X"01", --1688
  X"23", X"00", X"ED", X"B8", X"C1", X"78", X"0D", X"B9", --1690
  X"38", X"F4", X"EB", X"13", X"C1", X"E1", X"CD", X"2C", --1698
  X"36", X"01", X"23", X"00", X"ED", X"B0", X"37", X"C1", --16A0
  X"C9", X"E1", X"C1", X"C9", X"D5", X"26", X"00", X"68", --16A8
  X"19", X"57", X"78", X"5E", X"72", X"53", X"23", X"3C", --16B0
  X"FE", X"20", X"38", X"F7", X"7B", X"FE", X"00", X"D1", --16B8
  X"C9", X"D5", X"21", X"20", X"00", X"19", X"E5", X"57", --16C0
  X"3E", X"1F", X"18", X"07", X"5E", X"72", X"53", X"B8", --16C8
  X"28", X"04", X"3D", X"2B", X"18", X"F6", X"7B", X"FE", --16D0
  X"00", X"E1", X"D1", X"C9", X"B1", X"C9", X"BC", X"BE", --16D8
  X"C3", X"AF", X"B4", X"93", X"91", X"92", X"95", X"98", --16E0
  X"98", X"98", X"98", X"98", X"98", X"98", X"7F", X"81", --16E8
  X"2E", X"6C", X"6E", X"70", X"48", X"94", X"56", X"3F", --16F0
  X"41", X"2B", X"17", X"1F", X"37", X"77", X"44", X"0F", --16F8
  X"59", X"2B", X"43", X"2D", X"51", X"3A", X"6D", X"42", --1700
  X"0D", X"49", X"5C", X"44", X"15", X"5D", X"01", X"3D", --1708
  X"02", X"06", X"00", X"67", X"1E", X"06", X"CB", X"0E", --1710
  X"67", X"19", X"06", X"0C", X"53", X"1A", X"00", X"EE", --1718
  X"1C", X"0C", X"6F", X"1A", X"04", X"3D", X"06", X"CC", --1720
  X"06", X"0E", X"81", X"19", X"04", X"00", X"AB", X"1D", --1728
  X"0E", X"78", X"21", X"0E", X"8C", X"21", X"0E", X"D5", --1730
  X"21", X"0E", X"62", X"18", X"0C", X"AA", X"21", X"0D", --1738
  X"02", X"1A", X"0E", X"75", X"1B", X"08", X"00", X"80", --1740
  X"1E", X"03", X"4F", X"1E", X"00", X"5F", X"1E", X"0D", --1748
  X"0D", X"1A", X"00", X"6B", X"0D", X"09", X"00", X"DC", --1750
  X"22", X"06", X"00", X"3A", X"1F", X"0E", X"AB", X"19", --1758
  X"0E", X"EB", X"19", X"03", X"42", X"1E", X"09", X"0E", --1760
  X"BE", X"21", X"0C", X"A7", X"21", X"0E", X"74", X"21", --1768
  X"0E", X"71", X"1B", X"0B", X"0B", X"0B", X"0B", X"08", --1770
  X"00", X"F8", X"03", X"09", X"0E", X"AE", X"21", X"07", --1778
  X"07", X"07", X"07", X"07", X"07", X"08", X"00", X"7A", --1780
  X"1E", X"06", X"00", X"94", X"22", X"0E", X"8C", X"1A", --1788
  X"06", X"2C", X"0A", X"00", X"36", X"17", X"06", X"00", --1790
  X"E5", X"16", X"0E", X"41", X"06", X"0A", X"2C", X"0A", --1798
  X"0C", X"F0", X"1A", X"0E", X"0C", X"1C", X"0E", X"E5", --17A0
  X"1B", X"0C", X"2B", X"1B", X"0E", X"17", X"23", X"FD", --17A8
  X"CB", X"01", X"BE", X"EF", X"FB", X"19", X"AF", X"32", --17B0
  X"47", X"5C", X"3D", X"32", X"3A", X"5C", X"18", X"01", --17B8
  X"E7", X"EF", X"BF", X"16", X"FD", X"34", X"0D", X"FA", --17C0
  X"12", X"19", X"DF", X"06", X"00", X"FE", X"0D", X"CA", --17C8
  X"63", X"18", X"FE", X"3A", X"28", X"EA", X"21", X"21", --17D0
  X"18", X"E5", X"4F", X"E7", X"79", X"D6", X"CE", X"30", --17D8
  X"13", X"C6", X"CE", X"21", X"A9", X"17", X"FE", X"A3", --17E0
  X"28", X"16", X"21", X"AC", X"17", X"FE", X"A4", X"28", --17E8
  X"0F", X"C3", X"12", X"19", X"4F", X"21", X"DC", X"16", --17F0
  X"09", X"4E", X"09", X"18", X"03", X"2A", X"74", X"5C", --17F8
  X"7E", X"23", X"22", X"74", X"5C", X"01", X"FD", X"17", --1800
  X"C5", X"4F", X"FE", X"20", X"30", X"0C", X"21", X"B5", --1808
  X"18", X"06", X"00", X"09", X"4E", X"09", X"E5", X"DF", --1810
  X"05", X"C9", X"DF", X"B9", X"C2", X"12", X"19", X"E7", --1818
  X"C9", X"CD", X"D6", X"05", X"38", X"04", X"CD", X"AC", --1820
  X"05", X"14", X"FD", X"CB", X"0A", X"7E", X"C2", X"A8", --1828
  X"18", X"2A", X"42", X"5C", X"CB", X"7C", X"28", X"14", --1830
  X"21", X"FE", X"FF", X"22", X"45", X"5C", X"2A", X"61", --1838
  X"5C", X"2B", X"ED", X"5B", X"59", X"5C", X"1B", X"3A", --1840
  X"44", X"5C", X"18", X"36", X"EF", X"6E", X"19", X"3A", --1848
  X"44", X"5C", X"28", X"1C", X"A7", X"20", X"46", X"47", --1850
  X"7E", X"E6", X"C0", X"78", X"28", X"12", X"CD", X"AC", --1858
  X"05", X"FF", X"C1", X"FD", X"CB", X"01", X"7E", X"C8", --1860
  X"2A", X"55", X"5C", X"3E", X"C0", X"A6", X"C0", X"AF", --1868
  X"FE", X"01", X"CE", X"00", X"56", X"23", X"5E", X"ED", --1870
  X"53", X"45", X"5C", X"23", X"5E", X"23", X"56", X"EB", --1878
  X"19", X"23", X"22", X"55", X"5C", X"EB", X"22", X"5D", --1880
  X"5C", X"57", X"1E", X"00", X"FD", X"36", X"0A", X"FF", --1888
  X"15", X"FD", X"72", X"0D", X"CA", X"C0", X"17", X"14", --1890
  X"EF", X"8B", X"19", X"28", X"0B", X"CD", X"AC", X"05", --1898
  X"16", X"FD", X"CB", X"01", X"7E", X"C0", X"C1", X"C1", --18A0
  X"DF", X"FE", X"0D", X"28", X"B6", X"FE", X"3A", X"CA", --18A8
  X"C0", X"17", X"C3", X"12", X"19", X"24", X"43", X"46", --18B0
  X"1E", X"4C", X"20", X"53", X"5E", X"4D", X"86", X"57", --18B8
  X"88", X"06", X"02", X"05", X"EF", X"DE", X"1C", X"BF", --18C0
  X"C1", X"CC", X"A1", X"18", X"EB", X"2A", X"74", X"5C", --18C8
  X"4E", X"23", X"46", X"EB", X"C5", X"C9", X"EF", X"DE", --18D0
  X"1C", X"BF", X"C1", X"CC", X"A1", X"18", X"EB", X"2A", --18D8
  X"74", X"5C", X"4E", X"23", X"46", X"EB", X"E5", X"21", --18E0
  X"F8", X"18", X"22", X"5A", X"5B", X"21", X"14", X"5B", --18E8
  X"E3", X"E5", X"60", X"69", X"E3", X"C3", X"00", X"5B", --18F0
  X"C9", X"EF", X"1F", X"1C", X"C9", X"C1", X"EF", X"56", --18F8
  X"1C", X"CD", X"A1", X"18", X"C9", X"EF", X"6C", X"1C", --1900
  X"C9", X"E7", X"EF", X"7A", X"1C", X"C9", X"EF", X"82", --1908
  X"1C", X"C9", X"CD", X"AC", X"05", X"0B", X"EF", X"8C", --1910
  X"1C", X"C9", X"FD", X"CB", X"01", X"7E", X"FD", X"CB", --1918
  X"02", X"86", X"28", X"03", X"EF", X"4D", X"0D", X"F1", --1920
  X"3A", X"74", X"5C", X"D6", X"A7", X"EF", X"FC", X"21", --1928
  X"CD", X"A1", X"18", X"2A", X"8F", X"5C", X"22", X"8D", --1930
  X"5C", X"21", X"91", X"5C", X"7E", X"07", X"AE", X"E6", --1938
  X"AA", X"AE", X"77", X"C9", X"EF", X"BE", X"1C", X"C9", --1940
  X"F1", X"3A", X"66", X"5B", X"E6", X"0F", X"32", X"66", --1948
  X"5B", X"3A", X"74", X"5C", X"D6", X"74", X"32", X"74", --1950
  X"5C", X"CA", X"EB", X"11", X"3D", X"CA", X"F2", X"11", --1958
  X"3D", X"CA", X"F9", X"11", X"C3", X"00", X"12", X"C1", --1960
  X"FD", X"CB", X"01", X"7E", X"28", X"10", X"2A", X"65", --1968
  X"5C", X"11", X"FB", X"FF", X"19", X"22", X"65", X"5C", --1970
  X"EF", X"E9", X"34", X"DA", X"63", X"18", X"C3", X"C1", --1978
  X"17", X"FE", X"CD", X"20", X"09", X"E7", X"CD", X"0E", --1980
  X"19", X"CD", X"A1", X"18", X"18", X"18", X"CD", X"A1", --1988
  X"18", X"2A", X"65", X"5C", X"36", X"00", X"23", X"36", --1990
  X"00", X"23", X"36", X"01", X"23", X"36", X"00", X"23", --1998
  X"36", X"00", X"23", X"22", X"65", X"5C", X"EF", X"16", --19A0
  X"1D", X"C9", X"E7", X"CD", X"F9", X"18", X"FD", X"CB", --19A8
  X"01", X"7E", X"28", X"2E", X"DF", X"22", X"5F", X"5C", --19B0
  X"2A", X"57", X"5C", X"7E", X"FE", X"2C", X"28", X"0B", --19B8
  X"1E", X"E4", X"EF", X"86", X"1D", X"30", X"04", X"CD", --19C0
  X"AC", X"05", X"0D", X"23", X"22", X"5D", X"5C", X"7E", --19C8
  X"EF", X"56", X"1C", X"DF", X"22", X"57", X"5C", X"2A", --19D0
  X"5F", X"5C", X"FD", X"36", X"26", X"00", X"22", X"5D", --19D8
  X"5C", X"7E", X"DF", X"FE", X"2C", X"28", X"C3", X"CD", --19E0
  X"A1", X"18", X"C9", X"FD", X"CB", X"01", X"7E", X"20", --19E8
  X"0B", X"EF", X"FB", X"24", X"FE", X"2C", X"C4", X"A1", --19F0
  X"18", X"E7", X"18", X"F5", X"3E", X"E4", X"EF", X"39", --19F8
  X"1E", X"C9", X"EF", X"67", X"1E", X"01", X"00", X"00", --1A00
  X"EF", X"45", X"1E", X"18", X"03", X"EF", X"99", X"1E", --1A08
  X"78", X"B1", X"20", X"04", X"ED", X"4B", X"B2", X"5C", --1A10
  X"C5", X"ED", X"5B", X"4B", X"5C", X"2A", X"59", X"5C", --1A18
  X"2B", X"EF", X"E5", X"19", X"EF", X"6B", X"0D", X"2A", --1A20
  X"65", X"5C", X"11", X"32", X"00", X"19", X"D1", X"ED", --1A28
  X"52", X"30", X"08", X"2A", X"B4", X"5C", X"A7", X"ED", --1A30
  X"52", X"30", X"04", X"CD", X"AC", X"05", X"15", X"ED", --1A38
  X"53", X"B2", X"5C", X"D1", X"E1", X"C1", X"ED", X"7B", --1A40
  X"B2", X"5C", X"33", X"C5", X"E5", X"ED", X"73", X"3D", --1A48
  X"5C", X"D5", X"C9", X"D1", X"FD", X"66", X"0D", X"24", --1A50
  X"E3", X"33", X"ED", X"4B", X"45", X"5C", X"C5", X"E5", --1A58
  X"ED", X"73", X"3D", X"5C", X"D5", X"EF", X"67", X"1E", --1A60
  X"01", X"14", X"00", X"EF", X"05", X"1F", X"C9", X"C1", --1A68
  X"E1", X"D1", X"7A", X"FE", X"3E", X"28", X"0F", X"3B", --1A70
  X"E3", X"EB", X"ED", X"73", X"3D", X"5C", X"C5", X"22", --1A78
  X"42", X"5C", X"FD", X"72", X"0A", X"C9", X"D5", X"E5", --1A80
  X"CD", X"AC", X"05", X"06", X"FD", X"CB", X"01", X"7E", --1A88
  X"28", X"05", X"3E", X"CE", X"C3", X"FE", X"19", X"FD", --1A90
  X"CB", X"01", X"F6", X"EF", X"8D", X"2C", X"30", X"16", --1A98
  X"E7", X"FE", X"24", X"20", X"05", X"FD", X"CB", X"01", --1AA0
  X"B6", X"E7", X"FE", X"28", X"20", X"3C", X"E7", X"FE", --1AA8
  X"29", X"28", X"20", X"EF", X"8D", X"2C", X"D2", X"12", --1AB0
  X"19", X"EB", X"E7", X"FE", X"24", X"20", X"02", X"EB", --1AB8
  X"E7", X"EB", X"01", X"06", X"00", X"EF", X"55", X"16", --1AC0
  X"23", X"23", X"36", X"0E", X"FE", X"2C", X"20", X"03", --1AC8
  X"E7", X"18", X"E0", X"FE", X"29", X"20", X"13", X"E7", --1AD0
  X"FE", X"3D", X"20", X"0E", X"E7", X"3A", X"3B", X"5C", --1AD8
  X"F5", X"EF", X"FB", X"24", X"F1", X"FD", X"AE", X"01", --1AE0
  X"E6", X"40", X"C2", X"12", X"19", X"CD", X"A1", X"18", --1AE8
  X"C9", X"21", X"0E", X"EC", X"36", X"FF", X"CD", X"20", --1AF0
  X"1F", X"EF", X"B0", X"16", X"2A", X"59", X"5C", X"01", --1AF8
  X"03", X"00", X"EF", X"55", X"16", X"21", X"6E", X"1B", --1B00
  X"ED", X"5B", X"59", X"5C", X"01", X"03", X"00", X"ED", --1B08
  X"B0", X"CD", X"6B", X"02", X"CD", X"20", X"1F", X"EF", --1B10
  X"B0", X"16", X"2A", X"59", X"5C", X"01", X"01", X"00", --1B18
  X"EF", X"55", X"16", X"2A", X"59", X"5C", X"36", X"E1", --1B20
  X"CD", X"6B", X"02", X"CD", X"53", X"1B", X"ED", X"7B", --1B28
  X"3D", X"5C", X"E1", X"21", X"03", X"13", X"E5", X"21", --1B30
  X"13", X"00", X"E5", X"21", X"08", X"00", X"E5", X"3E", --1B38
  X"20", X"32", X"5C", X"5B", X"C3", X"00", X"5B", X"21", --1B40
  X"00", X"00", X"E5", X"3E", X"20", X"32", X"5C", X"5B", --1B48
  X"C3", X"00", X"5B", X"2A", X"4F", X"5C", X"11", X"05", --1B50
  X"00", X"19", X"11", X"0A", X"00", X"EB", X"19", X"EB", --1B58
  X"01", X"04", X"00", X"ED", X"B0", X"FD", X"CB", X"30", --1B60
  X"9E", X"FD", X"CB", X"01", X"A6", X"C9", X"EF", X"22", --1B68
  X"22", X"3E", X"03", X"18", X"02", X"3E", X"02", X"FD", --1B70
  X"36", X"02", X"00", X"EF", X"30", X"25", X"28", X"03", --1B78
  X"EF", X"01", X"16", X"EF", X"18", X"00", X"EF", X"70", --1B80
  X"20", X"38", X"18", X"EF", X"18", X"00", X"FE", X"3B", --1B88
  X"28", X"04", X"FE", X"2C", X"20", X"08", X"EF", X"20", --1B90
  X"00", X"CD", X"0E", X"19", X"18", X"08", X"EF", X"E6", --1B98
  X"1C", X"18", X"03", X"EF", X"DE", X"1C", X"CD", X"A1", --1BA0
  X"18", X"EF", X"25", X"18", X"C9", X"ED", X"73", X"81", --1BA8
  X"5B", X"31", X"FF", X"5B", X"CD", X"97", X"1C", X"ED", --1BB0
  X"4B", X"72", X"5B", X"21", X"F7", X"FF", X"F6", X"FF", --1BB8
  X"ED", X"42", X"CD", X"F3", X"1C", X"01", X"09", X"00", --1BC0
  X"21", X"71", X"5B", X"CD", X"AC", X"1D", X"2A", X"74", --1BC8
  X"5B", X"ED", X"4B", X"72", X"5B", X"CD", X"AC", X"1D", --1BD0
  X"CD", X"56", X"1D", X"3E", X"05", X"CD", X"64", X"1C", --1BD8
  X"ED", X"7B", X"81", X"5B", X"C9", X"EF", X"18", X"00", --1BE0
  X"FE", X"21", X"C2", X"12", X"19", X"EF", X"20", X"00", --1BE8
  X"CD", X"A1", X"18", X"3E", X"02", X"EF", X"01", X"16", --1BF0
  X"ED", X"73", X"81", X"5B", X"31", X"FF", X"5B", X"CD", --1BF8
  X"D2", X"20", X"3E", X"05", X"CD", X"64", X"1C", X"ED", --1C00
  X"7B", X"81", X"5B", X"C9", X"EF", X"18", X"00", X"FE", --1C08
  X"21", X"C2", X"12", X"19", X"CD", X"93", X"13", X"CD", --1C10
  X"A1", X"18", X"ED", X"73", X"81", X"5B", X"31", X"FF", --1C18
  X"5B", X"CD", X"5F", X"1F", X"3E", X"05", X"CD", X"64", --1C20
  X"1C", X"ED", X"7B", X"81", X"5B", X"C9", X"ED", X"73", --1C28
  X"81", X"5B", X"31", X"FF", X"5B", X"CD", X"35", X"1D", --1C30
  X"21", X"71", X"5B", X"01", X"09", X"00", X"CD", X"37", --1C38
  X"1E", X"3E", X"05", X"CD", X"64", X"1C", X"ED", X"7B", --1C40
  X"81", X"5B", X"C9", X"ED", X"73", X"81", X"5B", X"31", --1C48
  X"FF", X"5B", X"42", X"4B", X"CD", X"37", X"1E", X"CD", --1C50
  X"56", X"1D", X"3E", X"05", X"CD", X"64", X"1C", X"ED", --1C58
  X"7B", X"81", X"5B", X"C9", X"E5", X"C5", X"21", X"81", --1C60
  X"1C", X"06", X"00", X"4F", X"09", X"4E", X"F3", X"3A", --1C68
  X"5C", X"5B", X"E6", X"F8", X"B1", X"32", X"5C", X"5B", --1C70
  X"01", X"FD", X"7F", X"ED", X"79", X"FB", X"C1", X"E1", --1C78
  X"C9", X"01", X"03", X"04", X"06", X"07", X"00", X"11", --1C80
  X"67", X"5B", X"DD", X"E5", X"E1", X"06", X"0A", X"1A", --1C88
  X"13", X"BE", X"23", X"C0", X"10", X"F9", X"C9", X"CD", --1C90
  X"12", X"1D", X"28", X"04", X"CD", X"AC", X"05", X"20", --1C98
  X"DD", X"E5", X"01", X"EC", X"3F", X"DD", X"09", X"DD", --1CA0
  X"E1", X"30", X"63", X"21", X"EC", X"FF", X"3E", X"FF", --1CA8
  X"CD", X"F3", X"1C", X"21", X"66", X"5B", X"CB", X"D6", --1CB0
  X"DD", X"E5", X"D1", X"21", X"67", X"5B", X"01", X"0A", --1CB8
  X"00", X"ED", X"B0", X"DD", X"CB", X"13", X"C6", X"DD", --1CC0
  X"7E", X"0A", X"DD", X"77", X"10", X"DD", X"7E", X"0B", --1CC8
  X"DD", X"77", X"11", X"DD", X"7E", X"0C", X"DD", X"77", --1CD0
  X"12", X"AF", X"DD", X"77", X"0D", X"DD", X"77", X"0E", --1CD8
  X"DD", X"77", X"0F", X"3E", X"05", X"CD", X"64", X"1C", --1CE0
  X"DD", X"E5", X"E1", X"01", X"EC", X"FF", X"09", X"22", --1CE8
  X"83", X"5B", X"C9", X"ED", X"5B", X"85", X"5B", X"08", --1CF0
  X"3A", X"87", X"5B", X"4F", X"08", X"CB", X"7F", X"20", --1CF8
  X"09", X"19", X"89", X"22", X"85", X"5B", X"32", X"87", --1D00
  X"5B", X"C9", X"19", X"89", X"38", X"F5", X"CD", X"AC", --1D08
  X"05", X"03", X"3E", X"04", X"CD", X"64", X"1C", X"DD", --1D10
  X"21", X"EC", X"EB", X"ED", X"5B", X"83", X"5B", X"B7", --1D18
  X"DD", X"E5", X"E1", X"ED", X"52", X"C8", X"CD", X"87", --1D20
  X"1C", X"20", X"03", X"F6", X"FF", X"C9", X"01", X"EC", --1D28
  X"FF", X"DD", X"09", X"18", X"E6", X"CD", X"12", X"1D", --1D30
  X"20", X"04", X"CD", X"AC", X"05", X"23", X"DD", X"7E", --1D38
  X"0A", X"DD", X"77", X"10", X"DD", X"7E", X"0B", X"DD", --1D40
  X"77", X"11", X"DD", X"7E", X"0C", X"DD", X"77", X"12", --1D48
  X"3E", X"05", X"CD", X"64", X"1C", X"C9", X"3E", X"04", --1D50
  X"CD", X"64", X"1C", X"DD", X"CB", X"13", X"46", X"C8", --1D58
  X"DD", X"CB", X"13", X"86", X"21", X"66", X"5B", X"CB", --1D60
  X"96", X"DD", X"6E", X"10", X"DD", X"66", X"11", X"DD", --1D68
  X"7E", X"12", X"DD", X"5E", X"0A", X"DD", X"56", X"0B", --1D70
  X"DD", X"46", X"0C", X"B7", X"ED", X"52", X"98", X"CB", --1D78
  X"14", X"CB", X"14", X"CB", X"2F", X"CB", X"1C", X"CB", --1D80
  X"2F", X"CB", X"1C", X"DD", X"75", X"0D", X"DD", X"74", --1D88
  X"0E", X"DD", X"77", X"0F", X"DD", X"6E", X"10", X"DD", --1D90
  X"66", X"11", X"DD", X"7E", X"12", X"01", X"EC", X"FF", --1D98
  X"DD", X"09", X"DD", X"75", X"0A", X"DD", X"74", X"0B", --1DA0
  X"DD", X"77", X"0C", X"C9", X"78", X"B1", X"C8", X"E5", --1DA8
  X"11", X"00", X"C0", X"EB", X"ED", X"52", X"28", X"1D", --1DB0
  X"38", X"1B", X"E5", X"ED", X"42", X"30", X"0D", X"60", --1DB8
  X"69", X"C1", X"B7", X"ED", X"42", X"E3", X"11", X"00", --1DC0
  X"C0", X"D5", X"18", X"28", X"E1", X"E1", X"11", X"00", --1DC8
  X"00", X"D5", X"D5", X"18", X"1F", X"60", X"69", X"11", --1DD0
  X"20", X"00", X"B7", X"ED", X"52", X"38", X"05", X"E3", --1DD8
  X"42", X"4B", X"18", X"05", X"E1", X"11", X"00", X"00", --1DE0
  X"D5", X"C5", X"11", X"98", X"5B", X"ED", X"B0", X"C1", --1DE8
  X"E5", X"21", X"98", X"5B", X"3E", X"04", X"CD", X"64", --1DF0
  X"1C", X"DD", X"5E", X"10", X"DD", X"56", X"11", X"DD", --1DF8
  X"7E", X"12", X"CD", X"64", X"1C", X"ED", X"A0", X"7A", --1E00
  X"B3", X"28", X"19", X"78", X"B1", X"C2", X"05", X"1E", --1E08
  X"3E", X"04", X"CD", X"64", X"1C", X"DD", X"73", X"10", --1E10
  X"DD", X"72", X"11", X"3E", X"05", X"CD", X"64", X"1C", --1E18
  X"E1", X"C1", X"18", X"88", X"3E", X"04", X"CD", X"64", --1E20
  X"1C", X"DD", X"34", X"12", X"DD", X"7E", X"12", X"11", --1E28
  X"00", X"C0", X"CD", X"64", X"1C", X"18", X"D4", X"78", --1E30
  X"B1", X"C8", X"E5", X"11", X"00", X"C0", X"EB", X"ED", --1E38
  X"52", X"28", X"24", X"38", X"22", X"E5", X"ED", X"42", --1E40
  X"30", X"12", X"60", X"69", X"C1", X"B7", X"ED", X"42", --1E48
  X"E3", X"11", X"00", X"00", X"D5", X"11", X"00", X"C0", --1E50
  X"D5", X"EB", X"18", X"24", X"E1", X"E1", X"11", X"00", --1E58
  X"00", X"D5", X"D5", X"D5", X"EB", X"18", X"19", X"60", --1E60
  X"69", X"11", X"20", X"00", X"B7", X"ED", X"52", X"38", --1E68
  X"05", X"E3", X"42", X"4B", X"18", X"05", X"E1", X"11", --1E70
  X"00", X"00", X"D5", X"C5", X"E5", X"11", X"98", X"5B", --1E78
  X"3E", X"04", X"CD", X"64", X"1C", X"DD", X"6E", X"10", --1E80
  X"DD", X"66", X"11", X"DD", X"7E", X"12", X"CD", X"64", --1E88
  X"1C", X"ED", X"A0", X"7C", X"B5", X"28", X"25", X"78", --1E90
  X"B1", X"C2", X"91", X"1E", X"3E", X"04", X"CD", X"64", --1E98
  X"1C", X"DD", X"75", X"10", X"DD", X"74", X"11", X"3E", --1EA0
  X"05", X"CD", X"64", X"1C", X"D1", X"C1", X"21", X"98", --1EA8
  X"5B", X"78", X"B1", X"28", X"02", X"ED", X"B0", X"EB", --1EB0
  X"C1", X"C3", X"37", X"1E", X"3E", X"04", X"CD", X"64", --1EB8
  X"1C", X"DD", X"34", X"12", X"DD", X"7E", X"12", X"21", --1EC0
  X"00", X"C0", X"CD", X"64", X"1C", X"18", X"C8", X"F5", --1EC8
  X"3A", X"5C", X"5B", X"F5", X"E5", X"D5", X"C5", X"DD", --1ED0
  X"21", X"6A", X"5B", X"DD", X"73", X"10", X"DD", X"72", --1ED8
  X"11", X"DD", X"36", X"12", X"04", X"CD", X"AC", X"1D", --1EE0
  X"3E", X"05", X"CD", X"64", X"1C", X"C1", X"D1", X"E1", --1EE8
  X"09", X"EB", X"09", X"EB", X"F1", X"01", X"FD", X"7F", --1EF0
  X"F3", X"ED", X"79", X"32", X"5C", X"5B", X"FB", X"01", --1EF8
  X"00", X"00", X"F1", X"C9", X"F5", X"3A", X"5C", X"5B", --1F00
  X"F5", X"E5", X"D5", X"C5", X"DD", X"21", X"6A", X"5B", --1F08
  X"DD", X"75", X"10", X"DD", X"74", X"11", X"DD", X"36", --1F10
  X"12", X"04", X"EB", X"CD", X"37", X"1E", X"18", X"C8", --1F18
  X"08", X"3E", X"00", X"F3", X"CD", X"3A", X"1F", X"F1", --1F20
  X"22", X"58", X"5B", X"2A", X"81", X"5B", X"ED", X"73", --1F28
  X"81", X"5B", X"F9", X"FB", X"2A", X"58", X"5B", X"F5", --1F30
  X"08", X"C9", X"C5", X"01", X"FD", X"7F", X"ED", X"79", --1F38
  X"32", X"5C", X"5B", X"C1", X"C9", X"08", X"F3", X"F1", --1F40
  X"22", X"58", X"5B", X"2A", X"81", X"5B", X"ED", X"73", --1F48
  X"81", X"5B", X"F9", X"2A", X"58", X"5B", X"F5", X"3E", --1F50
  X"07", X"CD", X"3A", X"1F", X"FB", X"08", X"C9", X"CD", --1F58
  X"12", X"1D", X"20", X"04", X"CD", X"AC", X"05", X"23", --1F60
  X"DD", X"6E", X"0D", X"DD", X"66", X"0E", X"DD", X"7E", --1F68
  X"0F", X"CD", X"F3", X"1C", X"FD", X"E5", X"FD", X"2A", --1F70
  X"83", X"5B", X"01", X"EC", X"FF", X"DD", X"09", X"FD", --1F78
  X"6E", X"0A", X"FD", X"66", X"0B", X"FD", X"7E", X"0C", --1F80
  X"FD", X"E1", X"DD", X"5E", X"0A", X"DD", X"56", X"0B", --1F88
  X"DD", X"46", X"0C", X"B7", X"ED", X"52", X"98", X"CB", --1F90
  X"14", X"CB", X"14", X"CB", X"2F", X"CB", X"1C", X"CB", --1F98
  X"2F", X"CB", X"1C", X"01", X"14", X"00", X"DD", X"09", --1FA0
  X"DD", X"75", X"10", X"DD", X"74", X"11", X"DD", X"77", --1FA8
  X"12", X"01", X"EC", X"FF", X"DD", X"09", X"DD", X"6E", --1FB0
  X"0A", X"DD", X"66", X"0B", X"DD", X"56", X"0C", X"01", --1FB8
  X"14", X"00", X"DD", X"09", X"7A", X"CD", X"64", X"1C", --1FC0
  X"3A", X"5C", X"5B", X"5F", X"01", X"FD", X"7F", X"3E", --1FC8
  X"07", X"F3", X"ED", X"79", X"D9", X"DD", X"6E", X"0A", --1FD0
  X"DD", X"66", X"0B", X"DD", X"56", X"0C", X"7A", X"CD", --1FD8
  X"64", X"1C", X"3A", X"5C", X"5B", X"5F", X"01", X"FD", --1FE0
  X"7F", X"D9", X"3E", X"07", X"F3", X"ED", X"79", X"DD", --1FE8
  X"7E", X"10", X"D6", X"01", X"DD", X"77", X"10", X"30", --1FF0
  X"14", X"DD", X"7E", X"11", X"D6", X"01", X"DD", X"77", --1FF8
  X"11", X"30", X"0A", X"DD", X"7E", X"12", X"D6", X"01", --2000
  X"DD", X"77", X"12", X"38", X"31", X"ED", X"59", X"7E", --2008
  X"2C", X"20", X"11", X"24", X"20", X"0E", X"08", X"14", --2010
  X"7A", X"CD", X"64", X"1C", X"3A", X"5C", X"5B", X"5F", --2018
  X"21", X"00", X"C0", X"08", X"D9", X"F3", X"ED", X"59", --2020
  X"77", X"2C", X"20", X"0F", X"24", X"20", X"0C", X"14", --2028
  X"7A", X"CD", X"64", X"1C", X"3A", X"5C", X"5B", X"5F", --2030
  X"21", X"00", X"C0", X"D9", X"18", X"AC", X"3E", X"04", --2038
  X"CD", X"64", X"1C", X"3E", X"00", X"21", X"14", X"00", --2040
  X"CD", X"F3", X"1C", X"DD", X"5E", X"0D", X"DD", X"56", --2048
  X"0E", X"DD", X"4E", X"0F", X"7A", X"07", X"CB", X"11", --2050
  X"07", X"CB", X"11", X"7A", X"E6", X"3F", X"57", X"DD", --2058
  X"E5", X"D5", X"11", X"EC", X"FF", X"DD", X"19", X"D1", --2060
  X"DD", X"6E", X"0A", X"DD", X"66", X"0B", X"DD", X"7E", --2068
  X"0C", X"B7", X"ED", X"52", X"91", X"CB", X"74", X"20", --2070
  X"03", X"CB", X"F4", X"3D", X"DD", X"75", X"0A", X"DD", --2078
  X"74", X"0B", X"DD", X"77", X"0C", X"DD", X"6E", X"10", --2080
  X"DD", X"66", X"11", X"DD", X"7E", X"12", X"B7", X"ED", --2088
  X"52", X"91", X"CB", X"74", X"20", X"03", X"CB", X"F4", --2090
  X"3D", X"DD", X"75", X"10", X"DD", X"74", X"11", X"DD", --2098
  X"77", X"12", X"DD", X"E5", X"E1", X"D5", X"ED", X"5B", --20A0
  X"83", X"5B", X"B7", X"ED", X"52", X"D1", X"20", X"B1", --20A8
  X"ED", X"5B", X"83", X"5B", X"E1", X"E5", X"B7", X"ED", --20B0
  X"52", X"44", X"4D", X"E1", X"E5", X"11", X"14", X"00", --20B8
  X"19", X"EB", X"E1", X"1B", X"2B", X"ED", X"B8", X"2A", --20C0
  X"83", X"5B", X"11", X"14", X"00", X"19", X"22", X"83", --20C8
  X"5B", X"C9", X"3E", X"04", X"CD", X"64", X"1C", X"21", --20D0
  X"21", X"21", X"01", X"2B", X"21", X"DD", X"21", X"EC", --20D8
  X"EB", X"CD", X"D6", X"05", X"DD", X"E5", X"E3", X"ED", --20E0
  X"5B", X"83", X"5B", X"B7", X"ED", X"52", X"E1", X"28", --20E8
  X"20", X"54", X"5D", X"E5", X"C5", X"CD", X"8A", X"1C", --20F0
  X"C1", X"E1", X"30", X"0E", X"50", X"59", X"E5", X"C5", --20F8
  X"CD", X"8A", X"1C", X"C1", X"E1", X"38", X"03", X"DD", --2100
  X"E5", X"C1", X"11", X"EC", X"FF", X"DD", X"19", X"18", --2108
  X"D0", X"E5", X"21", X"2B", X"21", X"B7", X"ED", X"42", --2110
  X"E1", X"C8", X"60", X"69", X"CD", X"35", X"21", X"18", --2118
  X"B9", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --2120
  X"00", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"FF", --2128
  X"FF", X"FF", X"FF", X"FF", X"FF", X"E5", X"C5", X"E1", --2130
  X"11", X"67", X"5B", X"01", X"0A", X"00", X"ED", X"B0", --2138
  X"3E", X"05", X"CD", X"64", X"1C", X"2A", X"81", X"5B", --2140
  X"ED", X"73", X"81", X"5B", X"F9", X"21", X"67", X"5B", --2148
  X"06", X"0A", X"7E", X"E5", X"C5", X"EF", X"10", X"00", --2150
  X"C1", X"E1", X"23", X"10", X"F5", X"3E", X"0D", X"EF", --2158
  X"10", X"00", X"EF", X"4D", X"0D", X"2A", X"81", X"5B", --2160
  X"ED", X"73", X"81", X"5B", X"F9", X"3E", X"04", X"CD", --2168
  X"64", X"1C", X"E1", X"C9", X"3E", X"03", X"18", X"02", --2170
  X"3E", X"02", X"EF", X"30", X"25", X"28", X"03", X"EF", --2178
  X"01", X"16", X"EF", X"4D", X"0D", X"EF", X"DF", X"1F", --2180
  X"CD", X"A1", X"18", X"C9", X"EF", X"30", X"25", X"28", --2188
  X"08", X"3E", X"01", X"EF", X"01", X"16", X"EF", X"6E", --2190
  X"0D", X"FD", X"36", X"02", X"01", X"EF", X"C1", X"20", --2198
  X"CD", X"A1", X"18", X"EF", X"A0", X"20", X"C9", X"C3", --21A0
  X"F0", X"08", X"F3", X"C3", X"9D", X"01", X"DF", X"FE", --21A8
  X"2C", X"20", X"38", X"E7", X"EF", X"82", X"1C", X"CD", --21B0
  X"A1", X"18", X"EF", X"2D", X"23", X"C9", X"DF", X"FE", --21B8
  X"2C", X"28", X"07", X"CD", X"A1", X"18", X"EF", X"77", --21C0
  X"24", X"C9", X"E7", X"EF", X"82", X"1C", X"CD", X"A1", --21C8
  X"18", X"EF", X"94", X"23", X"C9", X"EF", X"B2", X"28", --21D0
  X"20", X"11", X"EF", X"30", X"25", X"20", X"08", X"CB", --21D8
  X"B1", X"EF", X"96", X"29", X"CD", X"A1", X"18", X"EF", --21E0
  X"15", X"2C", X"C9", X"CD", X"AC", X"05", X"0B", X"FD", --21E8
  X"CB", X"30", X"46", X"C8", X"EF", X"AF", X"0D", X"C9", --21F0
  X"21", X"FE", X"FF", X"22", X"45", X"5C", X"FD", X"CB", --21F8
  X"01", X"BE", X"CD", X"8E", X"22", X"EF", X"FB", X"24", --2200
  X"FD", X"CB", X"01", X"76", X"28", X"2C", X"DF", X"FE", --2208
  X"0D", X"20", X"27", X"FD", X"CB", X"01", X"FE", X"CD", --2210
  X"8E", X"22", X"21", X"21", X"03", X"22", X"8B", X"5B", --2218
  X"EF", X"FB", X"24", X"FD", X"CB", X"01", X"76", X"28", --2220
  X"11", X"11", X"8D", X"5B", X"2A", X"65", X"5C", X"01", --2228
  X"05", X"00", X"B7", X"ED", X"42", X"ED", X"B0", X"C3", --2230
  X"3E", X"22", X"CD", X"AC", X"05", X"19", X"3E", X"0D", --2238
  X"CD", X"6F", X"22", X"01", X"01", X"00", X"EF", X"30", --2240
  X"00", X"22", X"5B", X"5C", X"E5", X"2A", X"51", X"5C", --2248
  X"E5", X"3E", X"FF", X"EF", X"01", X"16", X"EF", X"E3", --2250
  X"2D", X"E1", X"EF", X"15", X"16", X"D1", X"2A", X"5B", --2258
  X"5C", X"A7", X"ED", X"52", X"1A", X"CD", X"6F", X"22", --2260
  X"13", X"2B", X"7C", X"B5", X"20", X"F6", X"C9", X"E5", --2268
  X"D5", X"CD", X"45", X"1F", X"21", X"0D", X"EC", X"CB", --2270
  X"9E", X"F5", X"3E", X"02", X"EF", X"01", X"16", X"F1", --2278
  X"CD", X"69", X"26", X"21", X"0D", X"EC", X"CB", X"9E", --2280
  X"CD", X"20", X"1F", X"D1", X"E1", X"C9", X"2A", X"59", --2288
  X"5C", X"2B", X"22", X"5D", X"5C", X"E7", X"C9", X"CD", --2290
  X"8E", X"22", X"FE", X"F1", X"C0", X"2A", X"5D", X"5C", --2298
  X"7E", X"23", X"FE", X"0D", X"C8", X"FE", X"3A", X"20", --22A0
  X"F7", X"B7", X"C9", X"47", X"21", X"BD", X"22", X"7E", --22A8
  X"23", X"B7", X"28", X"05", X"B8", X"20", X"F8", X"78", --22B0
  X"C9", X"F6", X"FF", X"78", X"C9", X"2B", X"2D", X"2A", --22B8
  X"2F", X"5E", X"3D", X"3E", X"3C", X"C7", X"C8", X"C9", --22C0
  X"C5", X"C6", X"00", X"FE", X"A5", X"38", X"0E", X"FE", --22C8
  X"C4", X"30", X"0A", X"FE", X"AC", X"28", X"06", X"FE", --22D0
  X"AD", X"28", X"02", X"BF", X"C9", X"FE", X"A5", X"C9", --22D8
  X"47", X"F6", X"20", X"FE", X"61", X"38", X"06", X"FE", --22E0
  X"7B", X"30", X"02", X"BF", X"C9", X"78", X"FE", X"2E", --22E8
  X"C8", X"CD", X"0A", X"23", X"20", X"11", X"E7", X"CD", --22F0
  X"0A", X"23", X"28", X"FA", X"FE", X"2E", X"C8", X"FE", --22F8
  X"45", X"C8", X"FE", X"65", X"C8", X"18", X"A4", X"F6", --2300
  X"FF", X"C9", X"FE", X"30", X"38", X"06", X"FE", X"3A", --2308
  X"30", X"02", X"BF", X"C9", X"FE", X"30", X"C9", X"06", --2310
  X"00", X"DF", X"C5", X"EF", X"8C", X"1C", X"C1", X"04", --2318
  X"FE", X"2C", X"20", X"03", X"E7", X"18", X"F3", X"78", --2320
  X"FE", X"09", X"38", X"04", X"CD", X"AC", X"05", X"2B", --2328
  X"CD", X"A1", X"18", X"C3", X"85", X"09", X"21", X"FF", --2330
  X"5B", X"22", X"81", X"5B", X"CD", X"45", X"1F", X"C3", --2338
  X"CB", X"25", X"A7", X"ED", X"52", X"44", X"4D", X"19", --2340
  X"EB", X"C9", X"01", X"01", X"00", X"E5", X"D5", X"CD", --2348
  X"58", X"23", X"D1", X"E1", X"EF", X"55", X"16", X"C9", --2350
  X"2A", X"65", X"5C", X"09", X"38", X"0A", X"EB", X"21", --2358
  X"82", X"00", X"19", X"38", X"03", X"ED", X"72", X"D8", --2360
  X"FD", X"36", X"00", X"03", X"C3", X"21", X"03", X"87", --2368
  X"87", X"6F", X"26", X"00", X"29", X"29", X"29", X"C9", --2370
  X"21", X"00", X"00", X"39", X"ED", X"5B", X"65", X"5C", --2378
  X"B7", X"ED", X"52", X"C9", X"FD", X"CB", X"C7", X"86", --2380
  X"CD", X"6F", X"23", X"E5", X"ED", X"5B", X"24", X"FF", --2388
  X"19", X"54", X"5D", X"E3", X"E5", X"D5", X"11", X"00", --2390
  X"58", X"19", X"EB", X"E1", X"01", X"20", X"00", X"3A", --2398
  X"8F", X"5C", X"CD", X"9B", X"24", X"E1", X"7C", X"26", --23A0
  X"00", X"87", X"87", X"87", X"C6", X"40", X"57", X"5C", --23A8
  X"19", X"EB", X"E1", X"06", X"20", X"C3", X"E1", X"23", --23B0
  X"16", X"FF", X"CD", X"6F", X"23", X"7A", X"ED", X"5B", --23B8
  X"24", X"FF", X"19", X"5D", X"54", X"13", X"77", X"0B", --23C0
  X"ED", X"B0", X"C9", X"CD", X"88", X"24", X"11", X"00", --23C8
  X"40", X"2A", X"24", X"FF", X"43", X"CD", X"E1", X"23", --23D0
  X"16", X"48", X"CD", X"E1", X"23", X"16", X"50", X"06", --23D8
  X"C0", X"7E", X"E5", X"D5", X"FE", X"FE", X"38", X"04", --23E0
  X"D6", X"FE", X"18", X"36", X"FE", X"20", X"30", X"07", --23E8
  X"21", X"27", X"25", X"A7", X"08", X"18", X"34", X"FE", --23F0
  X"80", X"30", X"0E", X"CD", X"71", X"23", X"ED", X"5B", --23F8
  X"36", X"5C", X"19", X"D1", X"CD", X"28", X"FF", X"18", --2400
  X"47", X"FE", X"90", X"30", X"04", X"D6", X"7F", X"18", --2408
  X"11", X"D6", X"90", X"CD", X"71", X"23", X"D1", X"CD", --2410
  X"20", X"1F", X"D5", X"ED", X"5B", X"7B", X"5C", X"37", --2418
  X"18", X"07", X"11", X"2F", X"25", X"CD", X"71", X"23", --2420
  X"A7", X"08", X"19", X"D1", X"4A", X"7E", X"12", X"23", --2428
  X"14", X"7E", X"12", X"23", X"14", X"7E", X"12", X"23", --2430
  X"14", X"7E", X"12", X"23", X"14", X"7E", X"12", X"23", --2438
  X"14", X"7E", X"12", X"23", X"14", X"7E", X"12", X"23", --2440
  X"14", X"7E", X"12", X"51", X"08", X"DC", X"45", X"1F", --2448
  X"E1", X"23", X"13", X"10", X"8C", X"C9", X"C5", X"F3", --2450
  X"01", X"FD", X"7F", X"3A", X"5C", X"5B", X"EE", X"10", --2458
  X"ED", X"79", X"FB", X"08", X"08", X"F3", X"0E", X"FD", --2460
  X"EE", X"10", X"ED", X"79", X"FB", X"C1", X"C9", X"21", --2468
  X"56", X"24", X"11", X"28", X"FF", X"01", X"0E", X"00", --2470
  X"ED", X"B0", X"E5", X"21", X"2C", X"24", X"0E", X"20", --2478
  X"ED", X"B0", X"E1", X"0E", X"0B", X"ED", X"B0", X"C9", --2480
  X"FD", X"CB", X"C7", X"86", X"11", X"00", X"58", X"01", --2488
  X"C0", X"02", X"2A", X"24", X"FF", X"3A", X"8D", X"5C", --2490
  X"32", X"8F", X"5C", X"08", X"C5", X"7E", X"FE", X"FF", --2498
  X"20", X"08", X"3A", X"8D", X"5C", X"12", X"23", X"13", --24A0
  X"18", X"5D", X"08", X"12", X"13", X"08", X"23", X"FE", --24A8
  X"15", X"30", X"54", X"FE", X"10", X"38", X"50", X"2B", --24B0
  X"20", X"08", X"23", X"7E", X"4F", X"08", X"E6", X"F8", --24B8
  X"18", X"43", X"FE", X"11", X"20", X"0B", X"23", X"7E", --24C0
  X"87", X"87", X"87", X"4F", X"08", X"E6", X"C7", X"18", --24C8
  X"34", X"FE", X"12", X"20", X"09", X"23", X"7E", X"0F", --24D0
  X"4F", X"08", X"E6", X"7F", X"18", X"27", X"FE", X"13", --24D8
  X"20", X"0A", X"23", X"7E", X"0F", X"0F", X"4F", X"08", --24E0
  X"E6", X"BF", X"18", X"19", X"FE", X"14", X"23", X"20", --24E8
  X"16", X"4E", X"3A", X"01", X"5C", X"A9", X"1F", X"30", --24F0
  X"0E", X"3E", X"01", X"FD", X"AE", X"C7", X"32", X"01", --24F8
  X"5C", X"08", X"CD", X"13", X"25", X"B1", X"08", X"C1", --2500
  X"0B", X"78", X"B1", X"C2", X"9C", X"24", X"08", X"32", --2508
  X"8F", X"5C", X"C9", X"47", X"E6", X"C0", X"4F", X"78", --2510
  X"87", X"87", X"87", X"E6", X"38", X"B1", X"4F", X"78", --2518
  X"1F", X"1F", X"1F", X"E6", X"07", X"B1", X"C9", X"00", --2520
  X"3C", X"62", X"60", X"6E", X"62", X"3E", X"00", X"00", --2528
  X"6C", X"10", X"54", X"BA", X"38", X"54", X"82", X"15", --2530
  X"0B", X"94", X"2A", X"0A", X"B5", X"2A", X"08", X"D7", --2538
  X"2A", X"09", X"E3", X"2A", X"AD", X"4F", X"2A", X"AC", --2540
  X"25", X"2A", X"AF", X"D4", X"29", X"AE", X"E1", X"29", --2548
  X"A6", X"83", X"29", X"A5", X"AB", X"29", X"A8", X"87", --2550
  X"2A", X"A7", X"7A", X"2A", X"AA", X"1B", X"29", X"0C", --2558
  X"2B", X"29", X"B3", X"17", X"30", X"B4", X"BC", X"2F", --2560
  X"B0", X"72", X"30", X"B1", X"3E", X"30", X"0D", X"44", --2568
  X"29", X"A9", X"9B", X"26", X"07", X"04", X"27", X"04", --2570
  X"0B", X"2E", X"27", X"0A", X"31", X"27", X"07", X"17", --2578
  X"27", X"0D", X"17", X"27", X"CD", X"BE", X"28", X"21", --2580
  X"00", X"00", X"22", X"9A", X"FC", X"3E", X"82", X"32", --2588
  X"0D", X"EC", X"21", X"00", X"00", X"22", X"49", X"5C", --2590
  X"CD", X"BC", X"35", X"CD", X"5E", X"36", X"C9", X"21", --2598
  X"FF", X"5B", X"22", X"81", X"5B", X"CD", X"45", X"1F", --25A0
  X"3E", X"02", X"EF", X"01", X"16", X"21", X"44", X"27", --25A8
  X"22", X"EA", X"F6", X"21", X"54", X"27", X"22", X"EC", --25B0
  X"F6", X"E5", X"21", X"0D", X"EC", X"CB", X"CE", X"CB", --25B8
  X"A6", X"2B", X"36", X"00", X"E1", X"CD", X"A8", X"36", --25C0
  X"C3", X"53", X"26", X"DD", X"21", X"6C", X"FD", X"21", --25C8
  X"FF", X"5B", X"22", X"81", X"5B", X"CD", X"45", X"1F", --25D0
  X"3E", X"02", X"EF", X"01", X"16", X"CD", X"68", X"36", --25D8
  X"21", X"3B", X"5C", X"CB", X"6E", X"28", X"FC", X"21", --25E0
  X"0D", X"EC", X"CB", X"9E", X"CB", X"76", X"20", X"14", --25E8
  X"3A", X"0E", X"EC", X"FE", X"04", X"28", X"0A", X"FE", --25F0
  X"00", X"C2", X"C7", X"28", X"CD", X"48", X"38", X"18", --25F8
  X"03", X"CD", X"4D", X"38", X"CD", X"D6", X"30", X"CD", --2600
  X"22", X"32", X"3A", X"0E", X"EC", X"FE", X"04", X"28", --2608
  X"42", X"2A", X"49", X"5C", X"7C", X"B5", X"20", X"15", --2610
  X"2A", X"53", X"5C", X"ED", X"4B", X"4B", X"5C", X"A7", --2618
  X"ED", X"42", X"20", X"06", X"21", X"00", X"00", X"22", --2620
  X"08", X"EC", X"2A", X"08", X"EC", X"CD", X"20", X"1F", --2628
  X"EF", X"6E", X"19", X"EF", X"95", X"16", X"CD", X"45", --2630
  X"1F", X"ED", X"53", X"49", X"5C", X"21", X"0D", X"EC", --2638
  X"CB", X"6E", X"20", X"0F", X"21", X"00", X"00", X"22", --2640
  X"06", X"EC", X"CD", X"2F", X"15", X"CD", X"F2", X"29", --2648
  X"CD", X"44", X"29", X"31", X"FF", X"5B", X"CD", X"68", --2650
  X"36", X"CD", X"7F", X"36", X"F5", X"3A", X"39", X"5C", --2658
  X"CD", X"EC", X"26", X"F1", X"CD", X"69", X"26", X"18", --2660
  X"EA", X"21", X"0D", X"EC", X"CB", X"4E", X"F5", X"21", --2668
  X"77", X"25", X"20", X"03", X"21", X"37", X"25", X"CD", --2670
  X"CE", X"3F", X"20", X"05", X"D4", X"E7", X"26", X"F1", --2678
  X"C9", X"F1", X"28", X"05", X"AF", X"32", X"41", X"5C", --2680
  X"C9", X"21", X"0D", X"EC", X"CB", X"46", X"28", X"04", --2688
  X"CD", X"E7", X"26", X"C9", X"FE", X"A3", X"30", X"BB", --2690
  X"C3", X"F1", X"28", X"3A", X"0E", X"EC", X"FE", X"04", --2698
  X"C8", X"CD", X"30", X"16", X"21", X"0D", X"EC", X"CB", --26A0
  X"9E", X"7E", X"EE", X"40", X"77", X"E6", X"40", X"28", --26A8
  X"05", X"CD", X"BB", X"26", X"18", X"03", X"CD", X"CE", --26B0
  X"26", X"37", X"C9", X"CD", X"81", X"38", X"21", X"0D", --26B8
  X"EC", X"CB", X"F6", X"CD", X"2D", X"2E", X"CD", X"88", --26C0
  X"3A", X"CD", X"DF", X"28", X"18", X"0B", X"21", X"0D", --26C8
  X"EC", X"CB", X"B6", X"CD", X"BE", X"28", X"CD", X"48", --26D0
  X"38", X"2A", X"9A", X"FC", X"7C", X"B5", X"C4", X"4A", --26D8
  X"33", X"CD", X"2F", X"15", X"C3", X"F2", X"29", X"3A", --26E0
  X"38", X"5C", X"CB", X"3F", X"DD", X"E5", X"16", X"00", --26E8
  X"5F", X"21", X"80", X"0C", X"EF", X"B5", X"03", X"DD", --26F0
  X"E1", X"C9", X"DD", X"E5", X"11", X"30", X"00", X"21", --26F8
  X"00", X"03", X"18", X"F0", X"CD", X"EC", X"29", X"21", --2700
  X"0D", X"EC", X"CB", X"CE", X"2B", X"36", X"00", X"2A", --2708
  X"EC", X"F6", X"CD", X"A8", X"36", X"37", X"C9", X"21", --2710
  X"0D", X"EC", X"CB", X"8E", X"2B", X"7E", X"2A", X"EA", --2718
  X"F6", X"E5", X"F5", X"CD", X"3E", X"37", X"F1", X"E1", --2720
  X"CD", X"CE", X"3F", X"C3", X"F2", X"29", X"37", X"18", --2728
  X"01", X"A7", X"21", X"0C", X"EC", X"7E", X"E5", X"2A", --2730
  X"EC", X"F6", X"DC", X"A7", X"37", X"D4", X"B6", X"37", --2738
  X"E1", X"77", X"37", X"C9", X"05", X"00", X"31", X"28", --2740
  X"01", X"6C", X"28", X"02", X"85", X"28", X"03", X"47", --2748
  X"1B", X"04", X"16", X"28", X"06", X"31", X"32", X"38", --2750
  X"20", X"20", X"20", X"20", X"20", X"FF", X"54", X"61", --2758
  X"70", X"65", X"20", X"4C", X"6F", X"61", X"64", X"65", --2760
  X"F2", X"31", X"32", X"38", X"20", X"42", X"41", X"53", --2768
  X"49", X"C3", X"43", X"61", X"6C", X"63", X"75", X"6C", --2770
  X"61", X"74", X"6F", X"F2", X"34", X"38", X"20", X"42", --2778
  X"41", X"53", X"49", X"C3", X"54", X"61", X"70", X"65", --2780
  X"20", X"54", X"65", X"73", X"74", X"65", X"F2", X"A0", --2788
  X"05", X"00", X"42", X"27", X"01", X"51", X"28", X"02", --2790
  X"11", X"28", X"03", X"62", X"28", X"04", X"1C", X"28", --2798
  X"06", X"4F", X"70", X"74", X"69", X"6F", X"6E", X"73", --27A0
  X"20", X"FF", X"31", X"32", X"38", X"20", X"42", X"41", --27A8
  X"53", X"49", X"C3", X"52", X"65", X"6E", X"75", X"6D", --27B0
  X"62", X"65", X"F2", X"53", X"63", X"72", X"65", X"65", --27B8
  X"EE", X"50", X"72", X"69", X"6E", X"F4", X"45", X"78", --27C0
  X"69", X"F4", X"A0", X"02", X"00", X"42", X"27", X"01", --27C8
  X"1C", X"28", X"03", X"4F", X"70", X"74", X"69", X"6F", --27D0
  X"6E", X"73", X"20", X"FF", X"43", X"61", X"6C", X"63", --27D8
  X"75", X"6C", X"61", X"74", X"6F", X"F2", X"45", X"78", --27E0
  X"69", X"F4", X"A0", X"16", X"01", X"00", X"10", X"00", --27E8
  X"11", X"07", X"13", X"00", X"54", X"6F", X"20", X"63", --27F0
  X"61", X"6E", X"63", X"65", X"6C", X"20", X"2D", X"20", --27F8
  X"70", X"72", X"65", X"73", X"73", X"20", X"42", X"52", --2800
  X"45", X"41", X"4B", X"20", X"74", X"77", X"69", X"63", --2808
  X"E5", X"CD", X"9B", X"26", X"18", X"5E", X"CD", X"57", --2810
  X"38", X"CD", X"E9", X"3B", X"21", X"0D", X"EC", X"CB", --2818
  X"B6", X"CD", X"BE", X"28", X"06", X"00", X"16", X"17", --2820
  X"CD", X"5E", X"3B", X"CD", X"20", X"1F", X"C3", X"9F", --2828
  X"25", X"CD", X"52", X"38", X"21", X"3C", X"5C", X"CB", --2830
  X"C6", X"11", X"EB", X"27", X"CD", X"7D", X"05", X"CB", --2838
  X"86", X"CB", X"F6", X"3E", X"07", X"32", X"0E", X"EC", --2840
  X"01", X"00", X"00", X"CD", X"2B", X"37", X"C3", X"F1", --2848
  X"1A", X"CD", X"88", X"38", X"D4", X"E7", X"26", X"21", --2850
  X"00", X"00", X"22", X"49", X"5C", X"22", X"08", X"EC", --2858
  X"18", X"03", X"CD", X"14", X"1B", X"21", X"0D", X"EC", --2860
  X"CB", X"76", X"20", X"08", X"21", X"3C", X"5C", X"CB", --2868
  X"86", X"CD", X"48", X"38", X"21", X"0D", X"EC", X"CB", --2870
  X"AE", X"CB", X"A6", X"3E", X"00", X"21", X"90", X"27", --2878
  X"11", X"A0", X"27", X"18", X"2C", X"21", X"0D", X"EC", --2880
  X"CB", X"EE", X"CB", X"E6", X"CB", X"B6", X"CD", X"BE", --2888
  X"28", X"CD", X"4D", X"38", X"3E", X"04", X"32", X"0E", --2890
  X"EC", X"21", X"00", X"00", X"22", X"49", X"5C", X"CD", --2898
  X"2F", X"15", X"01", X"00", X"00", X"78", X"CD", X"F8", --28A0
  X"29", X"3E", X"04", X"21", X"CB", X"27", X"11", X"D2", --28A8
  X"27", X"32", X"0E", X"EC", X"22", X"EA", X"F6", X"ED", --28B0
  X"53", X"EC", X"F6", X"C3", X"04", X"26", X"CD", X"1F", --28B8
  X"2E", X"CD", X"7F", X"3A", X"C3", X"E8", X"28", X"06", --28C0
  X"00", X"16", X"17", X"CD", X"5E", X"3B", X"C3", X"AD", --28C8
  X"25", X"06", X"00", X"00", X"00", X"04", X"10", X"14", --28D0
  X"06", X"00", X"00", X"00", X"00", X"01", X"01", X"21", --28D8
  X"D8", X"28", X"11", X"EE", X"F6", X"C3", X"BA", X"3F", --28E0
  X"21", X"D1", X"28", X"11", X"EE", X"F6", X"C3", X"BA", --28E8
  X"3F", X"21", X"0D", X"EC", X"B7", X"B7", X"CB", X"46", --28F0
  X"C2", X"F2", X"29", X"CB", X"BE", X"CB", X"DE", X"E5", --28F8
  X"F5", X"CD", X"EC", X"29", X"F1", X"F5", X"CD", X"81", --2900
  X"2E", X"F1", X"78", X"CD", X"78", X"2B", X"E1", X"CB", --2908
  X"FE", X"D2", X"F2", X"29", X"78", X"DA", X"F8", X"29", --2910
  X"C3", X"F2", X"29", X"21", X"0D", X"EC", X"CB", X"DE", --2918
  X"CD", X"EC", X"29", X"CD", X"12", X"2F", X"37", X"78", --2920
  X"C3", X"F8", X"29", X"21", X"0D", X"EC", X"CB", X"86", --2928
  X"CB", X"DE", X"CD", X"EC", X"29", X"CD", X"5B", X"2B", --2930
  X"3F", X"DA", X"F2", X"29", X"CD", X"12", X"2F", X"37", --2938
  X"78", X"C3", X"F8", X"29", X"CD", X"EC", X"29", X"F5", --2940
  X"CD", X"B4", X"30", X"C5", X"06", X"00", X"CD", X"41", --2948
  X"2E", X"C1", X"38", X"0A", X"21", X"20", X"00", X"19", --2950
  X"7E", X"2F", X"E6", X"09", X"28", X"1C", X"3A", X"0D", --2958
  X"EC", X"CB", X"5F", X"28", X"05", X"CD", X"8E", X"2C", --2960
  X"30", X"15", X"CD", X"4C", X"2C", X"CD", X"78", X"2B", --2968
  X"CD", X"CE", X"2E", X"06", X"00", X"F1", X"37", X"C3", --2970
  X"F8", X"29", X"F1", X"37", X"C3", X"F2", X"29", X"F1", --2978
  X"C3", X"F2", X"29", X"3A", X"0E", X"EC", X"FE", X"04", --2980
  X"C8", X"CD", X"EC", X"29", X"21", X"00", X"00", X"CD", --2988
  X"20", X"1F", X"EF", X"6E", X"19", X"EF", X"95", X"16", --2990
  X"CD", X"45", X"1F", X"ED", X"53", X"49", X"5C", X"3E", --2998
  X"0F", X"CD", X"96", X"3A", X"CD", X"2F", X"15", X"37", --29A0
  X"C3", X"F2", X"29", X"3A", X"0E", X"EC", X"FE", X"04", --29A8
  X"C8", X"CD", X"EC", X"29", X"21", X"0F", X"27", X"CD", --29B0
  X"20", X"1F", X"EF", X"6E", X"19", X"EB", X"EF", X"95", --29B8
  X"16", X"CD", X"45", X"1F", X"ED", X"53", X"49", X"5C", --29C0
  X"3E", X"0F", X"CD", X"96", X"3A", X"CD", X"2F", X"15", --29C8
  X"37", X"C3", X"F2", X"29", X"CD", X"EC", X"29", X"CD", --29D0
  X"EA", X"2B", X"D2", X"F2", X"29", X"78", X"C3", X"F8", --29D8
  X"29", X"CD", X"EC", X"29", X"CD", X"09", X"2C", X"30", --29E0
  X"09", X"78", X"18", X"0C", X"CD", X"07", X"2A", X"C3", --29E8
  X"4F", X"36", X"CD", X"07", X"2A", X"C3", X"40", X"36", --29F0
  X"CD", X"11", X"2A", X"F5", X"C5", X"3E", X"0F", X"CD", --29F8
  X"96", X"3A", X"C1", X"F1", X"C3", X"40", X"36", X"21", --2A00
  X"EE", X"F6", X"4E", X"23", X"46", X"23", X"7E", X"23", --2A08
  X"C9", X"21", X"EE", X"F6", X"71", X"23", X"70", X"23", --2A10
  X"77", X"C9", X"E5", X"CD", X"B4", X"30", X"26", X"00", --2A18
  X"68", X"19", X"7E", X"E1", X"C9", X"CD", X"EC", X"29", --2A20
  X"5F", X"16", X"0A", X"D5", X"CD", X"30", X"2B", X"D1", --2A28
  X"30", X"C0", X"7B", X"CD", X"11", X"2A", X"43", X"CD", --2A30
  X"F9", X"2A", X"30", X"06", X"15", X"20", X"EC", X"7B", --2A38
  X"38", X"B6", X"D5", X"CD", X"0B", X"2B", X"D1", X"43", --2A40
  X"CD", X"F9", X"2A", X"7B", X"B7", X"18", X"A9", X"CD", --2A48
  X"EC", X"29", X"5F", X"16", X"0A", X"D5", X"CD", X"0B", --2A50
  X"2B", X"D1", X"30", X"96", X"7B", X"CD", X"11", X"2A", --2A58
  X"43", X"CD", X"02", X"2B", X"30", X"07", X"15", X"20", --2A60
  X"EC", X"7B", X"DA", X"F8", X"29", X"F5", X"CD", X"30", --2A68
  X"2B", X"06", X"00", X"CD", X"D4", X"2B", X"F1", X"C3", --2A70
  X"F8", X"29", X"CD", X"EC", X"29", X"CD", X"4C", X"2C", --2A78
  X"D2", X"F2", X"29", X"78", X"C3", X"F8", X"29", X"CD", --2A80
  X"EC", X"29", X"CD", X"31", X"2C", X"D2", X"F2", X"29", --2A88
  X"78", X"C3", X"F8", X"29", X"CD", X"EC", X"29", X"5F", --2A90
  X"D5", X"CD", X"0B", X"2B", X"D1", X"D2", X"F2", X"29", --2A98
  X"43", X"CD", X"02", X"2B", X"7B", X"DA", X"F8", X"29", --2AA0
  X"F5", X"CD", X"30", X"2B", X"06", X"00", X"CD", X"F9", --2AA8
  X"2A", X"F1", X"C3", X"F8", X"29", X"CD", X"EC", X"29", --2AB0
  X"5F", X"D5", X"CD", X"30", X"2B", X"D1", X"D2", X"F2", --2AB8
  X"29", X"43", X"CD", X"02", X"2B", X"7B", X"DA", X"F8", --2AC0
  X"29", X"D5", X"CD", X"0B", X"2B", X"D1", X"43", X"CD", --2AC8
  X"F9", X"2A", X"7B", X"B7", X"C3", X"F8", X"29", X"CD", --2AD0
  X"EC", X"29", X"CD", X"5B", X"2B", X"DA", X"F8", X"29", --2AD8
  X"C3", X"F2", X"29", X"CD", X"EC", X"29", X"CD", X"78", --2AE0
  X"2B", X"DA", X"F8", X"29", X"F5", X"CD", X"0B", X"2B", --2AE8
  X"06", X"1F", X"CD", X"DF", X"2B", X"F1", X"C3", X"F8", --2AF0
  X"29", X"D5", X"CD", X"D4", X"2B", X"D4", X"DF", X"2B", --2AF8
  X"D1", X"C9", X"D5", X"CD", X"DF", X"2B", X"D4", X"D4", --2B00
  X"2B", X"D1", X"C9", X"CD", X"7C", X"2C", X"30", X"1F", --2B08
  X"C5", X"CD", X"B4", X"30", X"06", X"00", X"CD", X"41", --2B10
  X"2E", X"D4", X"80", X"2F", X"C1", X"21", X"F1", X"F6", --2B18
  X"7E", X"B9", X"38", X"09", X"C5", X"CD", X"6F", X"16", --2B20
  X"C1", X"D8", X"79", X"B7", X"C8", X"0D", X"37", X"C9", --2B28
  X"C5", X"CD", X"B4", X"30", X"06", X"00", X"CD", X"41", --2B30
  X"2E", X"C1", X"38", X"03", X"C3", X"80", X"2F", X"CD", --2B38
  X"68", X"2C", X"30", X"16", X"21", X"F1", X"F6", X"23", --2B40
  X"79", X"BE", X"38", X"0C", X"C5", X"E5", X"CD", X"39", --2B48
  X"16", X"E1", X"C1", X"D8", X"23", X"7E", X"B9", X"C8", --2B50
  X"0C", X"37", X"C9", X"57", X"05", X"FA", X"66", X"2B", --2B58
  X"58", X"CD", X"DF", X"2B", X"7B", X"D8", X"D5", X"CD", --2B60
  X"0B", X"2B", X"D1", X"7B", X"D0", X"06", X"1F", X"CD", --2B68
  X"DF", X"2B", X"78", X"D8", X"7A", X"06", X"00", X"C9", --2B70
  X"57", X"04", X"3E", X"1F", X"B8", X"38", X"06", X"58", --2B78
  X"CD", X"D4", X"2B", X"7B", X"D8", X"05", X"C5", X"E5", --2B80
  X"21", X"0D", X"EC", X"CB", X"7E", X"20", X"31", X"CD", --2B88
  X"B4", X"30", X"21", X"20", X"00", X"19", X"7E", X"CB", --2B90
  X"4F", X"20", X"25", X"CB", X"CE", X"CB", X"9E", X"21", --2B98
  X"23", X"00", X"19", X"EB", X"E1", X"C1", X"F5", X"CD", --2BA0
  X"30", X"2B", X"F1", X"CD", X"B4", X"30", X"21", X"23", --2BA8
  X"00", X"19", X"EB", X"CB", X"87", X"CB", X"DF", X"CD", --2BB0
  X"D3", X"2E", X"CD", X"F4", X"35", X"78", X"37", X"C9", --2BB8
  X"E1", X"C1", X"D5", X"CD", X"30", X"2B", X"D1", X"78", --2BC0
  X"D0", X"06", X"00", X"CD", X"D4", X"2B", X"78", X"D8", --2BC8
  X"7B", X"06", X"00", X"C9", X"D5", X"E5", X"CD", X"B4", --2BD0
  X"30", X"CD", X"41", X"2E", X"C3", X"65", X"2C", X"D5", --2BD8
  X"E5", X"CD", X"B4", X"30", X"CD", X"63", X"2E", X"C3", --2BE0
  X"65", X"2C", X"D5", X"E5", X"CD", X"5B", X"2B", X"30", --2BE8
  X"16", X"CD", X"1A", X"2A", X"FE", X"20", X"28", X"F4", --2BF0
  X"CD", X"5B", X"2B", X"30", X"0A", X"CD", X"1A", X"2A", --2BF8
  X"FE", X"20", X"20", X"F4", X"CD", X"78", X"2B", X"18", --2C00
  X"5C", X"D5", X"E5", X"CD", X"78", X"2B", X"30", X"1B", --2C08
  X"CD", X"1A", X"2A", X"FE", X"20", X"20", X"F4", X"CD", --2C10
  X"78", X"2B", X"30", X"0F", X"CD", X"41", X"2E", X"30", --2C18
  X"0A", X"CD", X"1A", X"2A", X"FE", X"20", X"28", X"EF", --2C20
  X"37", X"18", X"3A", X"D4", X"5B", X"2B", X"B7", X"18", --2C28
  X"34", X"D5", X"E5", X"CD", X"B4", X"30", X"21", X"20", --2C30
  X"00", X"19", X"CB", X"46", X"20", X"07", X"CD", X"0B", --2C38
  X"2B", X"38", X"F0", X"18", X"20", X"06", X"00", X"CD", --2C40
  X"D4", X"2B", X"18", X"19", X"D5", X"E5", X"CD", X"B4", --2C48
  X"30", X"21", X"20", X"00", X"19", X"CB", X"5E", X"20", --2C50
  X"07", X"CD", X"30", X"2B", X"38", X"F0", X"18", X"05", --2C58
  X"06", X"1F", X"CD", X"DF", X"2B", X"E1", X"D1", X"C9", --2C60
  X"3A", X"0D", X"EC", X"CB", X"5F", X"37", X"C8", X"CD", --2C68
  X"B4", X"30", X"21", X"20", X"00", X"19", X"CB", X"5E", --2C70
  X"37", X"C8", X"18", X"12", X"3A", X"0D", X"EC", X"CB", --2C78
  X"5F", X"37", X"C8", X"CD", X"B4", X"30", X"21", X"20", --2C80
  X"00", X"19", X"CB", X"46", X"37", X"C8", X"3E", X"02", --2C88
  X"CD", X"B4", X"30", X"21", X"20", X"00", X"19", X"CB", --2C90
  X"46", X"20", X"08", X"0D", X"F2", X"90", X"2C", X"0E", --2C98
  X"00", X"3E", X"01", X"21", X"00", X"EC", X"11", X"03", --2CA0
  X"EC", X"F6", X"80", X"77", X"12", X"23", X"13", X"3E", --2CA8
  X"00", X"77", X"12", X"23", X"13", X"79", X"77", X"12", --2CB0
  X"21", X"00", X"00", X"22", X"06", X"EC", X"CD", X"5F", --2CB8
  X"33", X"CD", X"67", X"3C", X"DD", X"E5", X"CD", X"20", --2CC0
  X"1F", X"CD", X"6B", X"02", X"CD", X"45", X"1F", X"DD", --2CC8
  X"E1", X"3A", X"3A", X"5C", X"3C", X"20", X"18", X"21", --2CD0
  X"0D", X"EC", X"CB", X"9E", X"CD", X"5E", X"36", X"3A", --2CD8
  X"0E", X"EC", X"FE", X"04", X"C4", X"2F", X"15", X"CD", --2CE0
  X"FA", X"26", X"CD", X"07", X"2A", X"37", X"C9", X"21", --2CE8
  X"00", X"EC", X"11", X"03", X"EC", X"1A", X"CB", X"BF", --2CF0
  X"77", X"23", X"13", X"1A", X"77", X"23", X"13", X"1A", --2CF8
  X"77", X"CD", X"63", X"3C", X"38", X"04", X"ED", X"4B", --2D00
  X"06", X"EC", X"2A", X"06", X"EC", X"B7", X"ED", X"42", --2D08
  X"F5", X"E5", X"CD", X"07", X"2A", X"E1", X"F1", X"38", --2D10
  X"11", X"28", X"2A", X"E5", X"78", X"CD", X"5B", X"2B", --2D18
  X"E1", X"30", X"22", X"2B", X"7C", X"B5", X"20", X"F3", --2D20
  X"18", X"1B", X"E5", X"21", X"0D", X"EC", X"CB", X"BE", --2D28
  X"E1", X"EB", X"21", X"00", X"00", X"B7", X"ED", X"52", --2D30
  X"E5", X"78", X"CD", X"78", X"2B", X"E1", X"30", X"05", --2D38
  X"2B", X"7C", X"B5", X"20", X"F3", X"21", X"0D", X"EC", --2D40
  X"CB", X"FE", X"CD", X"11", X"2A", X"3E", X"17", X"CD", --2D48
  X"96", X"3A", X"B7", X"C9", X"21", X"00", X"EC", X"CB", --2D50
  X"7E", X"28", X"07", X"2A", X"06", X"EC", X"23", X"22", --2D58
  X"06", X"EC", X"21", X"00", X"EC", X"7E", X"23", X"46", --2D60
  X"23", X"4E", X"E5", X"E6", X"0F", X"21", X"85", X"2D", --2D68
  X"CD", X"CE", X"3F", X"5D", X"E1", X"28", X"02", X"3E", --2D70
  X"0D", X"71", X"2B", X"70", X"2B", X"F5", X"7E", X"E6", --2D78
  X"F0", X"B3", X"77", X"F1", X"C9", X"03", X"02", X"AC", --2D80
  X"2D", X"04", X"E9", X"2D", X"01", X"8F", X"2D", X"CD", --2D88
  X"B7", X"32", X"CD", X"0E", X"2E", X"30", X"07", X"FE", --2D90
  X"00", X"28", X"F7", X"2E", X"01", X"C9", X"0C", X"06", --2D98
  X"00", X"2A", X"DB", X"F9", X"79", X"BE", X"38", X"E7", --2DA0
  X"06", X"00", X"0E", X"00", X"E5", X"21", X"EE", X"F6", --2DA8
  X"7E", X"B9", X"20", X"0A", X"23", X"7E", X"B8", X"20", --2DB0
  X"05", X"21", X"00", X"EC", X"CB", X"BE", X"E1", X"CD", --2DB8
  X"B4", X"30", X"CD", X"0E", X"2E", X"30", X"07", X"FE", --2DC0
  X"00", X"28", X"E1", X"2E", X"02", X"C9", X"21", X"20", --2DC8
  X"00", X"19", X"CB", X"5E", X"28", X"05", X"2E", X"08", --2DD0
  X"3E", X"0D", X"C9", X"21", X"F3", X"F6", X"0C", X"7E", --2DD8
  X"B9", X"06", X"00", X"30", X"DA", X"06", X"00", X"0E", --2DE0
  X"01", X"CD", X"C3", X"31", X"CD", X"0E", X"2E", X"30", --2DE8
  X"07", X"FE", X"00", X"28", X"F7", X"2E", X"04", X"C9", --2DF0
  X"21", X"20", X"00", X"19", X"CB", X"5E", X"20", X"09", --2DF8
  X"0C", X"06", X"00", X"3A", X"F5", X"F6", X"B9", X"30", --2E00
  X"E0", X"2E", X"08", X"3E", X"0D", X"C9", X"3E", X"1F", --2E08
  X"B8", X"3F", X"D0", X"68", X"26", X"00", X"19", X"7E", --2E10
  X"04", X"37", X"C9", X"01", X"14", X"01", X"01", X"21", --2E18
  X"3C", X"5C", X"CB", X"86", X"21", X"1B", X"2E", X"11", --2E20
  X"15", X"EC", X"C3", X"BA", X"3F", X"21", X"3C", X"5C", --2E28
  X"CB", X"C6", X"01", X"00", X"00", X"CD", X"2B", X"37", --2E30
  X"21", X"1D", X"2E", X"11", X"15", X"EC", X"C3", X"BA", --2E38
  X"3F", X"26", X"00", X"68", X"19", X"7E", X"FE", X"00", --2E40
  X"37", X"C0", X"78", X"B7", X"28", X"0D", X"E5", X"2B", --2E48
  X"7E", X"FE", X"00", X"37", X"E1", X"C0", X"7E", X"FE", --2E50
  X"00", X"37", X"C0", X"23", X"04", X"78", X"FE", X"1F", --2E58
  X"38", X"F4", X"C9", X"26", X"00", X"68", X"19", X"7E", --2E60
  X"FE", X"00", X"37", X"C0", X"7E", X"FE", X"00", X"20", --2E68
  X"07", X"78", X"B7", X"C8", X"2B", X"05", X"18", X"F4", --2E70
  X"04", X"37", X"C9", X"26", X"00", X"68", X"19", X"7E", --2E78
  X"C9", X"21", X"0D", X"EC", X"B7", X"CB", X"46", X"C0", --2E80
  X"C5", X"F5", X"CD", X"B4", X"30", X"F1", X"CD", X"AC", --2E88
  X"16", X"F5", X"EB", X"CD", X"04", X"36", X"EB", X"F1", --2E90
  X"3F", X"28", X"31", X"F5", X"06", X"00", X"0C", X"3A", --2E98
  X"15", X"EC", X"B9", X"38", X"23", X"7E", X"5F", X"E6", --2EA0
  X"D7", X"BE", X"77", X"7B", X"CB", X"CE", X"F5", X"CD", --2EA8
  X"B4", X"30", X"F1", X"28", X"0D", X"CB", X"87", X"CD", --2EB0
  X"D3", X"2E", X"30", X"10", X"CD", X"F4", X"35", X"F1", --2EB8
  X"18", X"CC", X"CD", X"41", X"2E", X"F1", X"18", X"C6", --2EC0
  X"F1", X"CD", X"6E", X"31", X"C1", X"C9", X"CD", X"B4", --2EC8
  X"30", X"3E", X"09", X"C5", X"D5", X"41", X"21", X"EF", --2ED0
  X"2E", X"4F", X"C5", X"CD", X"75", X"16", X"C1", X"79", --2ED8
  X"30", X"0A", X"48", X"CD", X"B4", X"30", X"21", X"20", --2EE0
  X"00", X"19", X"77", X"37", X"D1", X"C1", X"C9", X"00", --2EE8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --2EF0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --2EF8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --2F00
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"09", --2F08
  X"00", X"00", X"C5", X"CD", X"B4", X"30", X"C5", X"21", --2F10
  X"20", X"00", X"19", X"CB", X"4E", X"3E", X"00", X"28", --2F18
  X"10", X"0C", X"21", X"23", X"00", X"19", X"EB", X"3A", --2F20
  X"15", X"EC", X"B9", X"30", X"EA", X"0D", X"CD", X"C9", --2F28
  X"31", X"E1", X"E5", X"CD", X"B4", X"30", X"E1", X"47", --2F30
  X"79", X"BD", X"78", X"F5", X"20", X"03", X"44", X"18", --2F38
  X"09", X"F5", X"E5", X"06", X"00", X"CD", X"41", X"2E", --2F40
  X"E1", X"F1", X"E5", X"21", X"F4", X"F6", X"CB", X"C6", --2F48
  X"28", X"02", X"CB", X"86", X"CD", X"C1", X"16", X"F5", --2F50
  X"C5", X"D5", X"21", X"F4", X"F6", X"CB", X"46", X"20", --2F58
  X"0E", X"06", X"00", X"CD", X"D4", X"2B", X"38", X"07", --2F60
  X"CD", X"80", X"2F", X"D1", X"C1", X"18", X"05", X"E1", --2F68
  X"C1", X"CD", X"04", X"36", X"F1", X"0D", X"47", X"E1", --2F70
  X"F1", X"78", X"C2", X"32", X"2F", X"37", X"C1", X"C9", --2F78
  X"21", X"20", X"00", X"19", X"7E", X"CB", X"46", X"20", --2F80
  X"29", X"F5", X"C5", X"79", X"B7", X"20", X"15", X"C5", --2F88
  X"2A", X"9A", X"FC", X"CD", X"4A", X"33", X"22", X"9A", --2F90
  X"FC", X"3A", X"DB", X"F9", X"4F", X"0D", X"CD", X"B7", --2F98
  X"32", X"C1", X"18", X"04", X"0D", X"CD", X"B4", X"30", --2FA0
  X"C1", X"F1", X"21", X"20", X"00", X"19", X"CB", X"8E", --2FA8
  X"B6", X"77", X"41", X"CD", X"B4", X"30", X"CD", X"DF", --2FB0
  X"30", X"C3", X"48", X"16", X"CD", X"84", X"30", X"E5", --2FB8
  X"CD", X"95", X"30", X"28", X"32", X"CD", X"5B", X"2B", --2FC0
  X"E1", X"30", X"2D", X"CD", X"1A", X"2A", X"F5", X"E5", --2FC8
  X"CD", X"12", X"2F", X"E1", X"F1", X"FE", X"20", X"28", --2FD0
  X"E6", X"E5", X"CD", X"95", X"30", X"28", X"18", X"CD", --2FD8
  X"5B", X"2B", X"E1", X"30", X"13", X"CD", X"1A", X"2A", --2FE0
  X"FE", X"20", X"28", X"07", X"E5", X"CD", X"12", X"2F", --2FE8
  X"E1", X"18", X"E6", X"E5", X"CD", X"78", X"2B", X"E1", --2FF0
  X"78", X"F5", X"E5", X"21", X"F5", X"EE", X"CB", X"96", --2FF8
  X"3A", X"15", X"EC", X"C5", X"06", X"00", X"4F", X"BF", --3000
  X"CD", X"05", X"16", X"C1", X"21", X"0D", X"EC", X"CB", --3008
  X"DE", X"E1", X"CD", X"F8", X"29", X"F1", X"C9", X"CD", --3010
  X"84", X"30", X"E5", X"CD", X"1A", X"2A", X"E1", X"FE", --3018
  X"00", X"37", X"28", X"D4", X"F5", X"E5", X"CD", X"12", --3020
  X"2F", X"E1", X"F1", X"FE", X"20", X"20", X"EB", X"CD", --3028
  X"1A", X"2A", X"FE", X"20", X"37", X"20", X"C1", X"E5", --3030
  X"CD", X"12", X"2F", X"E1", X"18", X"F1", X"CD", X"84", --3038
  X"30", X"E5", X"CD", X"B4", X"30", X"21", X"20", X"00", --3040
  X"19", X"CB", X"46", X"20", X"0C", X"CD", X"5B", X"2B", --3048
  X"30", X"1B", X"CD", X"12", X"2F", X"E1", X"18", X"E9", --3050
  X"E5", X"78", X"FE", X"00", X"28", X"0F", X"05", X"CD", --3058
  X"1A", X"2A", X"04", X"FE", X"00", X"28", X"06", X"05", --3060
  X"CD", X"12", X"2F", X"18", X"EC", X"E1", X"37", X"C3", --3068
  X"F8", X"2F", X"CD", X"84", X"30", X"CD", X"1A", X"2A", --3070
  X"FE", X"00", X"37", X"28", X"F1", X"E5", X"CD", X"12", --3078
  X"2F", X"E1", X"18", X"F1", X"21", X"0D", X"EC", X"CB", --3080
  X"86", X"CD", X"EC", X"29", X"21", X"F5", X"EE", X"CB", --3088
  X"D6", X"21", X"F1", X"F6", X"C9", X"CD", X"B4", X"30", --3090
  X"21", X"20", X"00", X"19", X"CB", X"46", X"28", X"0E", --3098
  X"78", X"FE", X"00", X"28", X"0D", X"05", X"CD", X"1A", --30A0
  X"2A", X"04", X"FE", X"00", X"28", X"04", X"3E", X"01", --30A8
  X"B7", X"C9", X"AF", X"C9", X"21", X"16", X"EC", X"F5", --30B0
  X"79", X"11", X"23", X"00", X"B7", X"28", X"04", X"19", --30B8
  X"3D", X"18", X"F9", X"EB", X"F1", X"C9", X"D5", X"CD", --30C0
  X"B4", X"30", X"26", X"00", X"68", X"19", X"D1", X"C9", --30C8
  X"05", X"00", X"00", X"00", X"F8", X"F6", X"21", X"D0", --30D0
  X"30", X"11", X"F5", X"F6", X"C3", X"BA", X"3F", X"C5", --30D8
  X"D5", X"21", X"F5", X"F6", X"E5", X"7E", X"B7", X"20", --30E0
  X"18", X"E5", X"CD", X"5F", X"33", X"2A", X"D7", X"F9", --30E8
  X"CD", X"52", X"33", X"30", X"03", X"22", X"D7", X"F9", --30F0
  X"44", X"4D", X"E1", X"CD", X"D6", X"32", X"3D", X"18", --30F8
  X"15", X"21", X"0D", X"EC", X"CB", X"86", X"21", X"F8", --3100
  X"F6", X"54", X"5D", X"01", X"23", X"00", X"09", X"01", --3108
  X"BC", X"02", X"ED", X"B0", X"3D", X"37", X"D1", X"12", --3110
  X"21", X"F8", X"F6", X"D1", X"C1", X"C9", X"C5", X"D5", --3118
  X"21", X"20", X"00", X"19", X"7E", X"2F", X"E6", X"11", --3120
  X"20", X"15", X"E5", X"D5", X"23", X"56", X"23", X"5E", --3128
  X"D5", X"CD", X"5F", X"33", X"E1", X"CD", X"4A", X"33", --3130
  X"30", X"03", X"22", X"D7", X"F9", X"D1", X"E1", X"CB", --3138
  X"46", X"21", X"F5", X"F6", X"E5", X"28", X"05", X"3E", --3140
  X"00", X"37", X"18", X"CA", X"7E", X"FE", X"14", X"28", --3148
  X"C5", X"01", X"23", X"00", X"21", X"F8", X"F6", X"EB", --3150
  X"ED", X"B0", X"21", X"D6", X"F9", X"54", X"5D", X"01", --3158
  X"23", X"00", X"B7", X"ED", X"42", X"01", X"BC", X"02", --3160
  X"ED", X"B8", X"3C", X"37", X"18", X"A8", X"C5", X"D5", --3168
  X"F5", X"06", X"00", X"0E", X"01", X"E5", X"CD", X"C3", --3170
  X"31", X"E1", X"CB", X"5E", X"CB", X"9E", X"20", X"20", --3178
  X"CD", X"41", X"2E", X"F1", X"CD", X"AC", X"16", X"28", --3180
  X"31", X"F5", X"06", X"00", X"0C", X"79", X"FE", X"15", --3188
  X"38", X"0E", X"2B", X"7E", X"23", X"FE", X"00", X"28", --3190
  X"07", X"E5", X"21", X"0D", X"EC", X"CB", X"C6", X"E1", --3198
  X"CB", X"4E", X"CB", X"CE", X"CB", X"9E", X"CD", X"C3", --31A0
  X"31", X"20", X"D5", X"C5", X"D5", X"CD", X"E6", X"35", --31A8
  X"36", X"08", X"D1", X"C1", X"CD", X"F4", X"35", X"F1", --31B0
  X"18", X"CA", X"79", X"32", X"F5", X"F6", X"CB", X"DE", --31B8
  X"D1", X"C1", X"C9", X"21", X"F8", X"F6", X"C3", X"B7", --31C0
  X"30", X"C5", X"D5", X"21", X"0D", X"EC", X"CB", X"86", --31C8
  X"3A", X"F5", X"F6", X"4F", X"B7", X"3E", X"00", X"28", --31D0
  X"42", X"CD", X"C3", X"31", X"F5", X"06", X"00", X"CD", --31D8
  X"41", X"2E", X"30", X"0E", X"F1", X"CD", X"C1", X"16", --31E0
  X"F5", X"C5", X"06", X"00", X"CD", X"41", X"2E", X"C1", --31E8
  X"38", X"24", X"23", X"7E", X"F5", X"C5", X"79", X"FE", --31F0
  X"01", X"20", X"09", X"3A", X"15", X"EC", X"4F", X"CD", --31F8
  X"B4", X"30", X"18", X"04", X"0D", X"CD", X"C3", X"31", --3200
  X"C1", X"F1", X"21", X"20", X"00", X"19", X"CB", X"8E", --3208
  X"B6", X"77", X"21", X"F5", X"F6", X"35", X"F1", X"0D", --3210
  X"20", X"BF", X"37", X"D1", X"C1", X"C9", X"03", X"00", --3218
  X"DE", X"F9", X"21", X"1E", X"32", X"11", X"DB", X"F9", --3220
  X"C3", X"BA", X"3F", X"C5", X"D5", X"21", X"DB", X"F9", --3228
  X"E5", X"7E", X"B7", X"20", X"1E", X"E5", X"CD", X"5F", --3230
  X"33", X"2A", X"9A", X"FC", X"CD", X"4A", X"33", X"30", --3238
  X"03", X"22", X"9A", X"FC", X"44", X"4D", X"E1", X"23", --3240
  X"23", X"23", X"30", X"11", X"CD", X"D6", X"32", X"3D", --3248
  X"EB", X"18", X"0A", X"2A", X"DC", X"F9", X"01", X"23", --3250
  X"00", X"ED", X"42", X"37", X"3D", X"EB", X"E1", X"30", --3258
  X"01", X"77", X"23", X"73", X"23", X"72", X"EB", X"D1", --3260
  X"C1", X"C9", X"C5", X"D5", X"21", X"20", X"00", X"19", --3268
  X"7E", X"2F", X"E6", X"11", X"20", X"0C", X"D5", X"E5", --3270
  X"23", X"56", X"23", X"5E", X"ED", X"53", X"9A", X"FC", --3278
  X"E1", X"D1", X"CB", X"5E", X"21", X"DB", X"F9", X"E5", --3280
  X"28", X"16", X"E5", X"CD", X"5F", X"33", X"2A", X"9A", --3288
  X"FC", X"CD", X"52", X"33", X"22", X"9A", X"FC", X"E1", --3290
  X"23", X"23", X"23", X"3E", X"00", X"37", X"18", X"BD", --3298
  X"7E", X"FE", X"14", X"28", X"0E", X"3C", X"2A", X"DC", --32A0
  X"F9", X"01", X"23", X"00", X"EB", X"ED", X"B0", X"EB", --32A8
  X"37", X"18", X"AA", X"E1", X"D1", X"C1", X"C9", X"21", --32B0
  X"DE", X"F9", X"C3", X"B7", X"30", X"08", X"0D", X"CC", --32B8
  X"35", X"01", X"DA", X"35", X"12", X"5A", X"33", X"13", --32C0
  X"5A", X"33", X"14", X"5A", X"33", X"15", X"5A", X"33", --32C8
  X"10", X"5A", X"33", X"11", X"5A", X"33", X"54", X"5D", --32D0
  X"13", X"13", X"13", X"D5", X"21", X"20", X"00", X"19", --32D8
  X"36", X"01", X"23", X"70", X"23", X"71", X"0E", X"01", --32E0
  X"06", X"00", X"C5", X"D5", X"3A", X"0E", X"EC", X"FE", --32E8
  X"04", X"C4", X"17", X"35", X"D1", X"C1", X"38", X"0F", --32F0
  X"79", X"FE", X"01", X"3E", X"0D", X"20", X"08", X"78", --32F8
  X"B7", X"3E", X"01", X"28", X"02", X"3E", X"0D", X"21", --3300
  X"BD", X"32", X"CD", X"CE", X"3F", X"38", X"1D", X"28", --3308
  X"D9", X"F5", X"3E", X"1F", X"B8", X"30", X"0F", X"3E", --3310
  X"12", X"CD", X"31", X"33", X"38", X"05", X"F1", X"3E", --3318
  X"0D", X"18", X"E4", X"CD", X"F4", X"35", X"F1", X"CD", --3320
  X"C5", X"35", X"18", X"BE", X"E1", X"79", X"C8", X"37", --3328
  X"C9", X"F5", X"CD", X"E6", X"35", X"F1", X"AE", X"77", --3330
  X"79", X"FE", X"14", X"D0", X"0C", X"21", X"23", X"00", --3338
  X"19", X"EB", X"21", X"20", X"00", X"19", X"36", X"00", --3340
  X"37", X"C9", X"CD", X"B6", X"34", X"D8", X"21", X"00", --3348
  X"00", X"C9", X"CD", X"30", X"34", X"D8", X"21", X"00", --3350
  X"00", X"C9", X"CD", X"17", X"35", X"3F", X"D0", X"21", --3358
  X"00", X"00", X"22", X"9F", X"FC", X"22", X"A1", X"FC", --3360
  X"21", X"74", X"33", X"11", X"AE", X"FC", X"01", X"BC", --3368
  X"00", X"ED", X"B0", X"C9", X"F3", X"01", X"FD", X"7F", --3370
  X"16", X"17", X"ED", X"51", X"FE", X"50", X"30", X"31", --3378
  X"FE", X"40", X"30", X"26", X"FE", X"30", X"30", X"1B", --3380
  X"FE", X"20", X"30", X"10", X"FE", X"10", X"30", X"05", --3388
  X"21", X"96", X"00", X"18", X"21", X"D6", X"10", X"21", --3390
  X"CF", X"00", X"18", X"1A", X"D6", X"20", X"21", X"00", --3398
  X"01", X"18", X"13", X"D6", X"30", X"21", X"3E", X"01", --33A0
  X"18", X"0C", X"D6", X"40", X"21", X"8B", X"01", X"18", --33A8
  X"05", X"D6", X"50", X"21", X"D4", X"01", X"47", X"B7", --33B0
  X"28", X"09", X"7E", X"23", X"E6", X"80", X"28", X"FA", --33B8
  X"05", X"18", X"F5", X"11", X"A3", X"FC", X"ED", X"53", --33C0
  X"A1", X"FC", X"3A", X"9E", X"FC", X"B7", X"3E", X"00", --33C8
  X"32", X"9E", X"FC", X"20", X"04", X"3E", X"20", X"12", --33D0
  X"13", X"7E", X"47", X"23", X"12", X"13", X"E6", X"80", --33D8
  X"28", X"F7", X"78", X"E6", X"7F", X"1B", X"12", X"13", --33E0
  X"3E", X"A0", X"12", X"3E", X"07", X"01", X"FD", X"7F", --33E8
  X"ED", X"79", X"FB", X"C9", X"F3", X"01", X"FD", X"7F", --33F0
  X"16", X"17", X"ED", X"51", X"21", X"96", X"00", X"06", --33F8
  X"A5", X"11", X"74", X"FD", X"1A", X"E6", X"7F", X"FE", --3400
  X"61", X"1A", X"38", X"02", X"E6", X"DF", X"BE", X"20", --3408
  X"09", X"23", X"13", X"E6", X"80", X"28", X"ED", X"37", --3410
  X"18", X"0C", X"04", X"28", X"08", X"7E", X"E6", X"80", --3418
  X"23", X"28", X"FA", X"18", X"DC", X"B7", X"78", X"16", --3420
  X"07", X"01", X"FD", X"7F", X"ED", X"51", X"FB", X"C9", --3428
  X"CD", X"EA", X"34", X"B7", X"32", X"9E", X"FC", X"CD", --3430
  X"20", X"1F", X"CD", X"F6", X"34", X"30", X"52", X"20", --3438
  X"0C", X"78", X"B1", X"28", X"08", X"CD", X"CF", X"34", --3440
  X"CD", X"D9", X"34", X"30", X"44", X"56", X"23", X"5E", --3448
  X"CD", X"45", X"1F", X"D5", X"E5", X"DD", X"E5", X"DD", --3450
  X"21", X"A3", X"FC", X"DD", X"22", X"A1", X"FC", X"EB", --3458
  X"06", X"00", X"11", X"18", X"FC", X"CD", X"95", X"34", --3460
  X"11", X"9C", X"FF", X"CD", X"95", X"34", X"11", X"F6", --3468
  X"FF", X"CD", X"95", X"34", X"11", X"FF", X"FF", X"CD", --3470
  X"95", X"34", X"DD", X"2B", X"DD", X"7E", X"00", X"F6", --3478
  X"80", X"DD", X"77", X"00", X"DD", X"E1", X"E1", X"D1", --3480
  X"23", X"23", X"23", X"22", X"9F", X"FC", X"EB", X"37", --3488
  X"C9", X"CD", X"45", X"1F", X"C9", X"AF", X"19", X"3C", --3490
  X"38", X"FC", X"ED", X"52", X"3D", X"C6", X"30", X"DD", --3498
  X"77", X"00", X"FE", X"30", X"20", X"0B", X"78", X"B7", --34A0
  X"20", X"09", X"3E", X"00", X"DD", X"77", X"00", X"18", --34A8
  X"02", X"06", X"01", X"DD", X"23", X"C9", X"CD", X"EA", --34B0
  X"34", X"B7", X"32", X"9E", X"FC", X"CD", X"20", X"1F", --34B8
  X"CD", X"F6", X"34", X"30", X"CC", X"EB", X"7D", X"B4", --34C0
  X"37", X"C2", X"4D", X"34", X"3F", X"18", X"C2", X"E5", --34C8
  X"23", X"23", X"5E", X"23", X"56", X"23", X"19", X"D1", --34D0
  X"C9", X"7E", X"E6", X"C0", X"37", X"C8", X"3F", X"C9", --34D8
  X"78", X"BE", X"C0", X"79", X"23", X"BE", X"2B", X"C0", --34E0
  X"37", X"C9", X"E5", X"21", X"00", X"00", X"22", X"A1", --34E8
  X"FC", X"22", X"9F", X"FC", X"E1", X"C9", X"E5", X"C1", --34F0
  X"11", X"00", X"00", X"2A", X"53", X"5C", X"CD", X"D9", --34F8
  X"34", X"D0", X"CD", X"E0", X"34", X"D8", X"78", X"B1", --3500
  X"37", X"C8", X"CD", X"CF", X"34", X"CD", X"D9", X"34", --3508
  X"D0", X"CD", X"E0", X"34", X"30", X"F4", X"C9", X"2A", --3510
  X"A1", X"FC", X"7D", X"B4", X"28", X"1E", X"7E", X"23", --3518
  X"FE", X"A0", X"47", X"3E", X"00", X"20", X"02", X"3E", --3520
  X"FF", X"32", X"9E", X"FC", X"78", X"CB", X"7F", X"28", --3528
  X"03", X"21", X"00", X"00", X"22", X"A1", X"FC", X"E6", --3530
  X"7F", X"C3", X"8F", X"35", X"2A", X"9F", X"FC", X"7D", --3538
  X"B4", X"CA", X"91", X"35", X"CD", X"20", X"1F", X"7E", --3540
  X"FE", X"0E", X"20", X"08", X"23", X"23", X"23", X"23", --3548
  X"23", X"23", X"18", X"F3", X"CD", X"45", X"1F", X"23", --3550
  X"22", X"9F", X"FC", X"FE", X"A5", X"38", X"08", X"D6", --3558
  X"A5", X"CD", X"AE", X"FC", X"C3", X"17", X"35", X"FE", --3560
  X"A3", X"38", X"10", X"20", X"05", X"21", X"94", X"35", --3568
  X"18", X"03", X"21", X"9C", X"35", X"CD", X"FD", X"FC", --3570
  X"C3", X"17", X"35", X"F5", X"3E", X"00", X"32", X"9E", --3578
  X"FC", X"F1", X"FE", X"0D", X"20", X"09", X"21", X"00", --3580
  X"00", X"22", X"A1", X"FC", X"22", X"9F", X"FC", X"37", --3588
  X"C9", X"37", X"3F", X"C9", X"53", X"50", X"45", X"43", --3590
  X"54", X"52", X"55", X"CD", X"50", X"4C", X"41", X"D9", --3598
  X"47", X"4F", X"54", X"CF", X"47", X"4F", X"53", X"55", --35A0
  X"C2", X"44", X"45", X"46", X"46", X"CE", X"4F", X"50", --35A8
  X"45", X"4E", X"A3", X"43", X"4C", X"4F", X"53", X"45", --35B0
  X"A3", X"02", X"01", X"05", X"21", X"B9", X"35", X"11", --35B8
  X"6A", X"FD", X"C3", X"BA", X"3F", X"68", X"26", X"00", --35C0
  X"19", X"77", X"04", X"C9", X"CD", X"E6", X"35", X"7E", --35C8
  X"F6", X"18", X"77", X"21", X"6A", X"FD", X"CB", X"C6", --35D0
  X"37", X"C9", X"CD", X"E6", X"35", X"CB", X"DE", X"21", --35D8
  X"6A", X"FD", X"CB", X"C6", X"37", X"C9", X"68", X"26", --35E0
  X"00", X"19", X"3E", X"20", X"B8", X"C8", X"36", X"00", --35E8
  X"23", X"04", X"18", X"F8", X"3A", X"6B", X"FD", X"06", --35F0
  X"00", X"26", X"00", X"68", X"19", X"36", X"00", X"04", --35F8
  X"3D", X"20", X"F6", X"C9", X"C5", X"D5", X"E5", X"E5", --3600
  X"21", X"F5", X"EE", X"CB", X"56", X"E1", X"20", X"04", --3608
  X"41", X"CD", X"1E", X"3B", X"E1", X"D1", X"C1", X"C9", --3610
  X"C5", X"D5", X"E5", X"E5", X"21", X"F5", X"EE", X"CB", --3618
  X"56", X"E1", X"20", X"04", X"59", X"CD", X"BF", X"3A", --3620
  X"E1", X"D1", X"C1", X"C9", X"C5", X"D5", X"E5", X"E5", --3628
  X"21", X"F5", X"EE", X"CB", X"56", X"E1", X"20", X"04", --3630
  X"59", X"CD", X"C6", X"3A", X"E1", X"D1", X"C1", X"C9", --3638
  X"F5", X"C5", X"D5", X"E5", X"78", X"41", X"4F", X"CD", --3640
  X"9D", X"3A", X"E1", X"D1", X"C1", X"F1", X"C9", X"F5", --3648
  X"C5", X"D5", X"E5", X"78", X"41", X"4F", X"CD", X"B2", --3650
  X"3A", X"E1", X"D1", X"C1", X"F1", X"C9", X"3E", X"00", --3658
  X"32", X"41", X"5C", X"3E", X"02", X"32", X"0A", X"5C", --3660
  X"21", X"3B", X"5C", X"7E", X"F6", X"0C", X"77", X"21", --3668
  X"0D", X"EC", X"CB", X"66", X"21", X"66", X"5B", X"20", --3670
  X"03", X"CB", X"86", X"C9", X"CB", X"C6", X"C9", X"E5", --3678
  X"21", X"3B", X"5C", X"CB", X"6E", X"28", X"FC", X"CB", --3680
  X"AE", X"3A", X"08", X"5C", X"21", X"41", X"5C", X"CB", --3688
  X"86", X"FE", X"20", X"30", X"0D", X"FE", X"10", X"30", --3690
  X"E7", X"FE", X"06", X"38", X"E3", X"CD", X"A4", X"36", --3698
  X"30", X"DE", X"E1", X"C9", X"EF", X"DB", X"10", X"C9", --36A0
  X"E5", X"CD", X"3B", X"37", X"21", X"3C", X"5C", X"CB", --36A8
  X"86", X"E1", X"5E", X"23", X"E5", X"21", X"EC", X"37", --36B0
  X"CD", X"33", X"37", X"E1", X"CD", X"33", X"37", X"E5", --36B8
  X"CD", X"22", X"38", X"21", X"FA", X"37", X"CD", X"33", --36C0
  X"37", X"E1", X"D5", X"01", X"07", X"08", X"CD", X"2B", --36C8
  X"37", X"C5", X"06", X"0C", X"3E", X"20", X"D7", X"7E", --36D0
  X"23", X"FE", X"80", X"30", X"03", X"D7", X"10", X"F7", --36D8
  X"E6", X"7F", X"D7", X"3E", X"20", X"D7", X"10", X"FB", --36E0
  X"C1", X"04", X"CD", X"2B", X"37", X"1D", X"20", X"E1", --36E8
  X"21", X"38", X"6F", X"D1", X"CB", X"23", X"CB", X"23", --36F0
  X"CB", X"23", X"53", X"15", X"1E", X"6F", X"01", X"00", --36F8
  X"FF", X"7A", X"CD", X"19", X"37", X"01", X"01", X"00", --3700
  X"7B", X"CD", X"19", X"37", X"01", X"00", X"01", X"7A", --3708
  X"3C", X"CD", X"19", X"37", X"AF", X"CD", X"CA", X"37", --3710
  X"C9", X"F5", X"E5", X"D5", X"C5", X"44", X"4D", X"EF", --3718
  X"E9", X"22", X"C1", X"D1", X"E1", X"F1", X"09", X"3D", --3720
  X"20", X"EF", X"C9", X"3E", X"16", X"D7", X"78", X"D7", --3728
  X"79", X"D7", X"C9", X"7E", X"23", X"FE", X"FF", X"C8", --3730
  X"D7", X"18", X"F8", X"37", X"18", X"01", X"A7", X"11", --3738
  X"F6", X"EE", X"21", X"3C", X"5C", X"38", X"01", X"EB", --3740
  X"ED", X"A0", X"38", X"01", X"EB", X"21", X"7D", X"5C", --3748
  X"38", X"01", X"EB", X"01", X"14", X"00", X"ED", X"B0", --3750
  X"38", X"01", X"EB", X"08", X"01", X"07", X"07", X"CD", --3758
  X"94", X"3B", X"DD", X"7E", X"01", X"80", X"47", X"3E", --3760
  X"0C", X"C5", X"F5", X"D5", X"EF", X"9B", X"0E", X"01", --3768
  X"07", X"00", X"09", X"D1", X"CD", X"7E", X"37", X"F1", --3770
  X"C1", X"05", X"3D", X"20", X"EC", X"C9", X"01", X"0E", --3778
  X"08", X"C5", X"06", X"00", X"E5", X"08", X"38", X"01", --3780
  X"EB", X"ED", X"B0", X"38", X"01", X"EB", X"08", X"E1", --3788
  X"24", X"C1", X"10", X"ED", X"C5", X"D5", X"EF", X"88", --3790
  X"0E", X"EB", X"D1", X"C1", X"08", X"38", X"01", X"EB", --3798
  X"ED", X"B0", X"38", X"01", X"EB", X"08", X"C9", X"CD", --37A0
  X"CA", X"37", X"3D", X"F2", X"B1", X"37", X"7E", X"3D", --37A8
  X"3D", X"CD", X"CA", X"37", X"37", X"C9", X"D5", X"CD", --37B0
  X"CA", X"37", X"3C", X"57", X"7E", X"3D", X"3D", X"BA", --37B8
  X"7A", X"F2", X"C5", X"37", X"AF", X"CD", X"CA", X"37", --37C0
  X"D1", X"C9", X"F5", X"E5", X"D5", X"21", X"07", X"59", --37C8
  X"11", X"20", X"00", X"A7", X"28", X"04", X"19", X"3D", --37D0
  X"20", X"FC", X"3E", X"78", X"BE", X"20", X"02", X"3E", --37D8
  X"68", X"16", X"0E", X"77", X"23", X"15", X"20", X"FB", --37E0
  X"D1", X"E1", X"F1", X"C9", X"16", X"07", X"07", X"15", --37E8
  X"00", X"14", X"00", X"10", X"07", X"11", X"00", X"13", --37F0
  X"01", X"FF", X"11", X"00", X"20", X"11", X"07", X"10", --37F8
  X"00", X"FF", X"01", X"03", X"07", X"0F", X"1F", X"3F", --3800
  X"7F", X"FF", X"FE", X"FC", X"F8", X"F0", X"E0", X"C0", --3808
  X"80", X"00", X"10", X"02", X"20", X"11", X"06", X"21", --3810
  X"10", X"04", X"20", X"11", X"05", X"21", X"10", X"00", --3818
  X"20", X"FF", X"C5", X"D5", X"E5", X"21", X"02", X"38", --3820
  X"11", X"98", X"5B", X"01", X"10", X"00", X"ED", X"B0", --3828
  X"2A", X"36", X"5C", X"E5", X"21", X"98", X"5A", X"22", --3830
  X"36", X"5C", X"21", X"12", X"38", X"CD", X"33", X"37", --3838
  X"E1", X"22", X"36", X"5C", X"E1", X"D1", X"C1", X"C9", --3840
  X"21", X"69", X"27", X"18", X"0D", X"21", X"72", X"27", --3848
  X"18", X"08", X"21", X"5E", X"27", X"18", X"03", X"21", --3850
  X"84", X"27", X"E5", X"CD", X"81", X"38", X"21", X"A0", --3858
  X"5A", X"06", X"20", X"3E", X"40", X"77", X"23", X"10", --3860
  X"FC", X"21", X"EC", X"37", X"CD", X"33", X"37", X"01", --3868
  X"00", X"15", X"CD", X"2B", X"37", X"D1", X"CD", X"7D", --3870
  X"05", X"0E", X"1A", X"CD", X"2B", X"37", X"C3", X"22", --3878
  X"38", X"06", X"15", X"16", X"17", X"C3", X"5E", X"3B", --3880
  X"CD", X"20", X"1F", X"CD", X"05", X"3A", X"7A", X"B3", --3888
  X"CA", X"C0", X"39", X"2A", X"96", X"5B", X"EF", X"A9", --3890
  X"30", X"EB", X"2A", X"94", X"5B", X"19", X"11", X"10", --3898
  X"27", X"B7", X"ED", X"52", X"D2", X"C0", X"39", X"2A", --38A0
  X"53", X"5C", X"EF", X"B8", X"19", X"23", X"23", X"22", --38A8
  X"92", X"5B", X"23", X"23", X"ED", X"53", X"6B", X"5B", --38B0
  X"7E", X"EF", X"B6", X"18", X"FE", X"0D", X"28", X"05", --38B8
  X"CD", X"0E", X"39", X"18", X"F3", X"ED", X"5B", X"6B", --38C0
  X"5B", X"2A", X"4B", X"5C", X"A7", X"ED", X"52", X"EB", --38C8
  X"20", X"D8", X"CD", X"05", X"3A", X"42", X"4B", X"11", --38D0
  X"00", X"00", X"2A", X"53", X"5C", X"C5", X"D5", X"E5", --38D8
  X"2A", X"96", X"5B", X"EF", X"A9", X"30", X"ED", X"5B", --38E0
  X"94", X"5B", X"19", X"EB", X"E1", X"72", X"23", X"73", --38E8
  X"23", X"4E", X"23", X"46", X"23", X"09", X"D1", X"13", --38F0
  X"C1", X"0B", X"78", X"B1", X"20", X"DF", X"CD", X"45", --38F8
  X"1F", X"ED", X"43", X"92", X"5B", X"37", X"C9", X"CA", --3900
  X"F0", X"E1", X"EC", X"ED", X"E5", X"F7", X"23", X"22", --3908
  X"79", X"5B", X"EB", X"01", X"07", X"00", X"21", X"07", --3910
  X"39", X"ED", X"B1", X"EB", X"C0", X"0E", X"00", X"7E", --3918
  X"FE", X"20", X"28", X"1B", X"EF", X"1B", X"2D", X"30", --3920
  X"16", X"FE", X"2E", X"28", X"12", X"FE", X"0E", X"28", --3928
  X"12", X"F6", X"20", X"FE", X"65", X"20", X"04", X"78", --3930
  X"B1", X"20", X"04", X"2A", X"79", X"5B", X"C9", X"03", --3938
  X"23", X"18", X"DC", X"ED", X"43", X"71", X"5B", X"E5", --3940
  X"EF", X"B6", X"18", X"CD", X"36", X"3A", X"7E", X"E1", --3948
  X"FE", X"3A", X"28", X"03", X"FE", X"0D", X"C0", X"23", --3950
  X"EF", X"B4", X"33", X"EF", X"A2", X"2D", X"60", X"69", --3958
  X"EF", X"6E", X"19", X"28", X"0A", X"7E", X"FE", X"80", --3960
  X"20", X"05", X"21", X"0F", X"27", X"18", X"11", X"22", --3968
  X"77", X"5B", X"CD", X"0B", X"3A", X"2A", X"96", X"5B", --3970
  X"EF", X"A9", X"30", X"ED", X"5B", X"94", X"5B", X"19", --3978
  X"11", X"73", X"5B", X"E5", X"CD", X"3C", X"3A", X"58", --3980
  X"1C", X"16", X"00", X"D5", X"E5", X"6B", X"26", X"00", --3988
  X"ED", X"4B", X"71", X"5B", X"B7", X"ED", X"42", X"22", --3990
  X"71", X"5B", X"28", X"33", X"38", X"27", X"44", X"4D", --3998
  X"2A", X"79", X"5B", X"E5", X"D5", X"2A", X"65", X"5C", --39A0
  X"09", X"38", X"13", X"EB", X"21", X"82", X"00", X"19", --39A8
  X"38", X"0C", X"ED", X"72", X"3F", X"38", X"07", X"D1", --39B0
  X"E1", X"EF", X"55", X"16", X"18", X"11", X"D1", X"E1", --39B8
  X"CD", X"45", X"1F", X"A7", X"C9", X"0B", X"1D", X"20", --39C0
  X"FC", X"2A", X"79", X"5B", X"EF", X"E8", X"19", X"ED", --39C8
  X"5B", X"79", X"5B", X"E1", X"C1", X"ED", X"B0", X"EB", --39D0
  X"36", X"0E", X"C1", X"23", X"E5", X"EF", X"2B", X"2D", --39D8
  X"D1", X"01", X"05", X"00", X"ED", X"B0", X"EB", X"E5", --39E0
  X"2A", X"92", X"5B", X"E5", X"5E", X"23", X"56", X"2A", --39E8
  X"71", X"5B", X"19", X"EB", X"E1", X"73", X"23", X"72", --39F0
  X"2A", X"6B", X"5B", X"ED", X"5B", X"71", X"5B", X"19", --39F8
  X"22", X"6B", X"5B", X"E1", X"C9", X"2A", X"4B", X"5C", --3A00
  X"22", X"77", X"5B", X"2A", X"53", X"5C", X"ED", X"5B", --3A08
  X"77", X"5B", X"B7", X"ED", X"52", X"28", X"1A", X"2A", --3A10
  X"53", X"5C", X"01", X"00", X"00", X"C5", X"EF", X"B8", --3A18
  X"19", X"2A", X"77", X"5B", X"A7", X"ED", X"52", X"28", --3A20
  X"05", X"EB", X"C1", X"03", X"18", X"EF", X"D1", X"13", --3A28
  X"C9", X"11", X"00", X"00", X"C9", X"23", X"7E", X"FE", --3A30
  X"20", X"28", X"FA", X"C9", X"D5", X"01", X"18", X"FC", --3A38
  X"CD", X"60", X"3A", X"01", X"9C", X"FF", X"CD", X"60", --3A40
  X"3A", X"0E", X"F6", X"CD", X"60", X"3A", X"7D", X"C6", --3A48
  X"30", X"12", X"13", X"06", X"03", X"E1", X"7E", X"FE", --3A50
  X"30", X"C0", X"36", X"20", X"23", X"10", X"F7", X"C9", --3A58
  X"AF", X"09", X"3C", X"38", X"FC", X"ED", X"42", X"3D", --3A60
  X"C6", X"30", X"12", X"13", X"C9", X"08", X"00", X"00", --3A68
  X"14", X"00", X"00", X"00", X"0F", X"00", X"08", X"00", --3A70
  X"16", X"01", X"00", X"00", X"00", X"0F", X"00", X"DD", --3A78
  X"21", X"6C", X"FD", X"21", X"6D", X"3A", X"18", X"03", --3A80
  X"21", X"76", X"3A", X"11", X"6C", X"FD", X"C3", X"BA", --3A88
  X"3F", X"D7", X"7A", X"D7", X"37", X"C9", X"E6", X"3F", --3A90
  X"DD", X"77", X"06", X"37", X"C9", X"DD", X"7E", X"01", --3A98
  X"80", X"47", X"CD", X"A0", X"3B", X"7E", X"DD", X"77", --3AA0
  X"07", X"2F", X"E6", X"C0", X"DD", X"B6", X"06", X"77", --3AA8
  X"37", X"C9", X"DD", X"7E", X"01", X"80", X"47", X"CD", --3AB0
  X"A0", X"3B", X"DD", X"7E", X"07", X"77", X"C9", X"E5", --3AB8
  X"26", X"00", X"7B", X"90", X"18", X"07", X"E5", X"7B", --3AC0
  X"58", X"47", X"93", X"26", X"FF", X"4F", X"78", X"BB", --3AC8
  X"28", X"4B", X"D5", X"CD", X"98", X"3B", X"C5", X"4C", --3AD0
  X"EF", X"9B", X"0E", X"EB", X"AF", X"B1", X"28", X"03", --3AD8
  X"04", X"18", X"01", X"05", X"D5", X"EF", X"9B", X"0E", --3AE0
  X"D1", X"79", X"0E", X"20", X"06", X"08", X"C5", X"E5", --3AE8
  X"D5", X"06", X"00", X"ED", X"B0", X"D1", X"E1", X"C1", --3AF0
  X"24", X"14", X"10", X"F2", X"F5", X"D5", X"EF", X"88", --3AF8
  X"0E", X"EB", X"E3", X"EF", X"88", X"0E", X"EB", X"E3", --3B00
  X"D1", X"01", X"20", X"00", X"ED", X"B0", X"F1", X"C1", --3B08
  X"A7", X"28", X"03", X"04", X"18", X"01", X"05", X"0D", --3B10
  X"67", X"20", X"BB", X"D1", X"43", X"E1", X"CD", X"B8", --3B18
  X"3B", X"EB", X"3A", X"3C", X"5C", X"F5", X"21", X"0D", --3B20
  X"EC", X"CB", X"76", X"CB", X"87", X"28", X"02", X"CB", --3B28
  X"C7", X"32", X"3C", X"5C", X"0E", X"00", X"CD", X"2B", --3B30
  X"37", X"EB", X"06", X"20", X"7E", X"A7", X"20", X"02", --3B38
  X"3E", X"20", X"FE", X"90", X"30", X"0F", X"EF", X"10", --3B40
  X"00", X"23", X"10", X"F0", X"F1", X"32", X"3C", X"5C", --3B48
  X"CD", X"B8", X"3B", X"37", X"C9", X"CD", X"20", X"1F", --3B50
  X"D7", X"CD", X"45", X"1F", X"18", X"EB", X"CD", X"B8", --3B58
  X"3B", X"7A", X"90", X"3C", X"4F", X"CD", X"98", X"3B", --3B60
  X"C5", X"EF", X"9B", X"0E", X"0E", X"08", X"E5", X"06", --3B68
  X"20", X"AF", X"77", X"23", X"10", X"FC", X"E1", X"24", --3B70
  X"0D", X"20", X"F3", X"06", X"20", X"C5", X"EF", X"88", --3B78
  X"0E", X"EB", X"C1", X"3A", X"8D", X"5C", X"77", X"23", --3B80
  X"10", X"FC", X"C1", X"05", X"0D", X"20", X"D9", X"CD", --3B88
  X"B8", X"3B", X"37", X"C9", X"3E", X"21", X"91", X"4F", --3B90
  X"3E", X"18", X"90", X"DD", X"96", X"01", X"47", X"C9", --3B98
  X"C5", X"AF", X"50", X"5F", X"CB", X"1A", X"CB", X"1B", --3BA0
  X"CB", X"1A", X"CB", X"1B", X"CB", X"1A", X"CB", X"1B", --3BA8
  X"21", X"00", X"58", X"47", X"09", X"19", X"C1", X"C9", --3BB0
  X"F5", X"E5", X"D5", X"2A", X"8D", X"5C", X"ED", X"5B", --3BB8
  X"8F", X"5C", X"D9", X"2A", X"0F", X"EC", X"ED", X"5B", --3BC0
  X"11", X"EC", X"22", X"8D", X"5C", X"ED", X"53", X"8F", --3BC8
  X"5C", X"D9", X"22", X"0F", X"EC", X"ED", X"53", X"11", --3BD0
  X"EC", X"21", X"13", X"EC", X"3A", X"91", X"5C", X"56", --3BD8
  X"77", X"7A", X"32", X"91", X"5C", X"D1", X"E1", X"F1", --3BE0
  X"C9", X"CD", X"56", X"3C", X"F3", X"DB", X"FE", X"E6", --3BE8
  X"40", X"08", X"21", X"E1", X"58", X"11", X"06", X"00", --3BF0
  X"43", X"7A", X"77", X"19", X"10", X"FC", X"21", X"00", --3BF8
  X"00", X"11", X"00", X"08", X"01", X"FE", X"BF", X"ED", --3C00
  X"78", X"CB", X"47", X"28", X"49", X"06", X"7F", X"ED", --3C08
  X"78", X"CB", X"47", X"28", X"41", X"06", X"F7", X"ED", --3C10
  X"78", X"CB", X"47", X"28", X"39", X"1B", X"7A", X"B3", --3C18
  X"28", X"09", X"DB", X"FE", X"E6", X"40", X"28", X"F5", --3C20
  X"23", X"18", X"F2", X"CB", X"15", X"CB", X"14", X"CB", --3C28
  X"15", X"CB", X"14", X"08", X"28", X"07", X"08", X"3E", --3C30
  X"20", X"94", X"6F", X"18", X"02", X"08", X"6C", X"AF", --3C38
  X"67", X"11", X"1F", X"59", X"06", X"20", X"3E", X"48", --3C40
  X"FB", X"76", X"F3", X"12", X"1B", X"10", X"FC", X"13", --3C48
  X"19", X"3E", X"68", X"77", X"18", X"A8", X"FB", X"06", --3C50
  X"19", X"76", X"10", X"FD", X"21", X"3B", X"5C", X"CB", --3C58
  X"AE", X"37", X"C9", X"3E", X"01", X"18", X"02", X"3E", --3C60
  X"00", X"32", X"8A", X"FD", X"21", X"00", X"00", X"22", --3C68
  X"85", X"FD", X"22", X"87", X"FD", X"39", X"22", X"8B", --3C70
  X"FD", X"CD", X"EA", X"34", X"3E", X"00", X"32", X"84", --3C78
  X"FD", X"21", X"74", X"FD", X"22", X"7D", X"FD", X"CD", --3C80
  X"20", X"1F", X"EF", X"B0", X"16", X"CD", X"45", X"1F", --3C88
  X"3E", X"00", X"32", X"81", X"FD", X"2A", X"59", X"5C", --3C90
  X"22", X"82", X"FD", X"21", X"00", X"00", X"22", X"7F", --3C98
  X"FD", X"2A", X"85", X"FD", X"23", X"22", X"85", X"FD", --3CA0
  X"CD", X"9D", X"3D", X"4F", X"3A", X"81", X"FD", X"FE", --3CA8
  X"00", X"20", X"41", X"79", X"E6", X"04", X"28", X"35", --3CB0
  X"CD", X"E9", X"3D", X"30", X"07", X"3E", X"01", X"32", --3CB8
  X"81", X"FD", X"18", X"DD", X"2A", X"7F", X"FD", X"7D", --3CC0
  X"B4", X"C2", X"1E", X"3D", X"C5", X"CD", X"CD", X"3D", --3CC8
  X"C1", X"3E", X"00", X"32", X"81", X"FD", X"79", X"E6", --3CD0
  X"01", X"20", X"D8", X"78", X"CD", X"16", X"3E", X"D0", --3CD8
  X"2A", X"85", X"FD", X"23", X"22", X"85", X"FD", X"CD", --3CE0
  X"9D", X"3D", X"4F", X"18", X"E9", X"78", X"CD", X"16", --3CE8
  X"3E", X"D0", X"18", X"AD", X"FE", X"01", X"20", X"F5", --3CF0
  X"79", X"E6", X"01", X"28", X"BB", X"C5", X"CD", X"7E", --3CF8
  X"3F", X"C1", X"38", X"79", X"2A", X"7F", X"FD", X"7C", --3D00
  X"B5", X"20", X"13", X"79", X"E6", X"02", X"28", X"BC", --3D08
  X"CD", X"E9", X"3D", X"30", X"AF", X"2A", X"7D", X"FD", --3D10
  X"2B", X"22", X"7F", X"FD", X"18", X"83", X"C5", X"21", --3D18
  X"74", X"FD", X"ED", X"5B", X"7F", X"FD", X"7A", X"BC", --3D20
  X"20", X"05", X"7B", X"BD", X"20", X"01", X"13", X"1B", --3D28
  X"18", X"01", X"23", X"7E", X"E6", X"7F", X"E5", X"D5", --3D30
  X"CD", X"16", X"3E", X"D1", X"E1", X"7C", X"BA", X"20", --3D38
  X"F1", X"7D", X"BB", X"20", X"ED", X"ED", X"5B", X"7F", --3D40
  X"FD", X"21", X"74", X"FD", X"22", X"7F", X"FD", X"ED", --3D48
  X"4B", X"7D", X"FD", X"0B", X"7A", X"BC", X"20", X"18", --3D50
  X"7B", X"BD", X"20", X"14", X"13", X"E5", X"21", X"00", --3D58
  X"00", X"22", X"7F", X"FD", X"E1", X"78", X"BC", X"20", --3D60
  X"07", X"79", X"BD", X"20", X"03", X"C1", X"18", X"1F", --3D68
  X"1A", X"77", X"23", X"13", X"E6", X"80", X"28", X"F8", --3D70
  X"22", X"7D", X"FD", X"18", X"81", X"C5", X"CD", X"16", --3D78
  X"3E", X"C1", X"21", X"00", X"00", X"22", X"7F", X"FD", --3D80
  X"3A", X"81", X"FD", X"FE", X"04", X"28", X"05", X"3E", --3D88
  X"00", X"32", X"81", X"FD", X"21", X"74", X"FD", X"22", --3D90
  X"7D", X"FD", X"C3", X"B3", X"3C", X"CD", X"54", X"2D", --3D98
  X"47", X"FE", X"3F", X"38", X"0A", X"F6", X"20", X"CD", --3DA0
  X"C6", X"3D", X"38", X"17", X"3E", X"01", X"C9", X"FE", --3DA8
  X"20", X"28", X"0D", X"FE", X"23", X"28", X"06", X"38", --3DB0
  X"F3", X"FE", X"24", X"20", X"EF", X"3E", X"02", X"C9", --3DB8
  X"3E", X"03", X"C9", X"3E", X"06", X"C9", X"FE", X"7B", --3DC0
  X"D0", X"FE", X"61", X"3F", X"C9", X"21", X"74", X"FD", --3DC8
  X"22", X"7D", X"FD", X"97", X"32", X"7F", X"FD", X"32", --3DD0
  X"80", X"FD", X"7E", X"E6", X"7F", X"E5", X"CD", X"9C", --3DD8
  X"3E", X"E1", X"7E", X"E6", X"80", X"C0", X"23", X"18", --3DE0
  X"F1", X"2A", X"7D", X"FD", X"11", X"7D", X"FD", X"7A", --3DE8
  X"BC", X"20", X"05", X"7B", X"BD", X"CA", X"13", X"3E", --3DF0
  X"11", X"74", X"FD", X"7A", X"BC", X"20", X"04", X"7B", --3DF8
  X"BD", X"28", X"06", X"2B", X"7E", X"E6", X"7F", X"77", --3E00
  X"23", X"78", X"F6", X"80", X"77", X"23", X"22", X"7D", --3E08
  X"FD", X"37", X"C9", X"37", X"3F", X"C9", X"F5", X"3A", --3E10
  X"89", X"FD", X"B7", X"20", X"12", X"F1", X"FE", X"3E", --3E18
  X"28", X"08", X"FE", X"3C", X"28", X"04", X"CD", X"64", --3E20
  X"3E", X"C9", X"32", X"89", X"FD", X"37", X"C9", X"FE", --3E28
  X"3C", X"3E", X"00", X"32", X"89", X"FD", X"20", X"1A", --3E30
  X"F1", X"FE", X"3E", X"20", X"04", X"3E", X"C9", X"18", --3E38
  X"E5", X"FE", X"3D", X"20", X"04", X"3E", X"C7", X"18", --3E40
  X"DD", X"F5", X"3E", X"3C", X"CD", X"64", X"3E", X"F1", --3E48
  X"18", X"D4", X"F1", X"FE", X"3D", X"20", X"04", X"3E", --3E50
  X"C8", X"18", X"CB", X"F5", X"3E", X"3E", X"CD", X"64", --3E58
  X"3E", X"F1", X"18", X"C2", X"FE", X"0D", X"28", X"20", --3E60
  X"FE", X"EA", X"47", X"20", X"07", X"3E", X"04", X"32", --3E68
  X"81", X"FD", X"18", X"0E", X"FE", X"22", X"20", X"0A", --3E70
  X"3A", X"81", X"FD", X"E6", X"FE", X"EE", X"02", X"32", --3E78
  X"81", X"FD", X"78", X"CD", X"9C", X"3E", X"37", X"C9", --3E80
  X"3A", X"8A", X"FD", X"FE", X"00", X"28", X"0A", X"ED", --3E88
  X"4B", X"85", X"FD", X"2A", X"8B", X"FD", X"F9", X"37", --3E90
  X"C9", X"37", X"3F", X"C9", X"5F", X"3A", X"84", X"FD", --3E98
  X"57", X"7B", X"FE", X"20", X"20", X"20", X"7A", X"E6", --3EA0
  X"01", X"20", X"14", X"7A", X"E6", X"02", X"20", X"07", --3EA8
  X"7A", X"F6", X"02", X"32", X"84", X"FD", X"C9", X"7B", --3EB0
  X"CD", X"FB", X"3E", X"3A", X"84", X"FD", X"C9", X"7A", --3EB8
  X"E6", X"FE", X"32", X"84", X"FD", X"C9", X"FE", X"A3", --3EC0
  X"30", X"24", X"7A", X"E6", X"02", X"20", X"0B", X"7A", --3EC8
  X"E6", X"FE", X"32", X"84", X"FD", X"7B", X"CD", X"FB", --3ED0
  X"3E", X"C9", X"D5", X"3E", X"20", X"CD", X"FB", X"3E", --3ED8
  X"D1", X"7A", X"E6", X"FE", X"E6", X"FD", X"32", X"84", --3EE0
  X"FD", X"7B", X"CD", X"FB", X"3E", X"C9", X"7A", X"E6", --3EE8
  X"FD", X"F6", X"01", X"32", X"84", X"FD", X"7B", X"CD", --3EF0
  X"FB", X"3E", X"C9", X"2A", X"87", X"FD", X"23", X"22", --3EF8
  X"87", X"FD", X"2A", X"82", X"FD", X"47", X"3A", X"8A", --3F00
  X"FD", X"FE", X"00", X"78", X"28", X"25", X"ED", X"5B", --3F08
  X"5F", X"5C", X"7C", X"BA", X"20", X"1A", X"7D", X"BB", --3F10
  X"20", X"16", X"ED", X"4B", X"85", X"FD", X"2A", X"87", --3F18
  X"FD", X"A7", X"ED", X"42", X"30", X"04", X"ED", X"4B", --3F20
  X"87", X"FD", X"2A", X"8B", X"FD", X"F9", X"37", X"C9", --3F28
  X"37", X"18", X"02", X"37", X"3F", X"CD", X"20", X"1F", --3F30
  X"30", X"0D", X"7E", X"EB", X"FE", X"0E", X"20", X"1D", --3F38
  X"13", X"13", X"13", X"13", X"13", X"18", X"16", X"F5", --3F40
  X"01", X"01", X"00", X"E5", X"D5", X"CD", X"66", X"3F", --3F48
  X"D1", X"E1", X"EF", X"64", X"16", X"2A", X"65", X"5C", --3F50
  X"EB", X"ED", X"B8", X"F1", X"12", X"13", X"CD", X"45", --3F58
  X"1F", X"ED", X"53", X"82", X"FD", X"C9", X"2A", X"65", --3F60
  X"5C", X"09", X"38", X"0A", X"EB", X"21", X"82", X"00", --3F68
  X"19", X"38", X"03", X"ED", X"72", X"D8", X"3E", X"03", --3F70
  X"32", X"3A", X"5C", X"C3", X"21", X"03", X"CD", X"2E", --3F78
  X"FD", X"D8", X"06", X"F9", X"11", X"74", X"FD", X"21", --3F80
  X"94", X"35", X"CD", X"3B", X"FD", X"D0", X"FE", X"FF", --3F88
  X"20", X"04", X"3E", X"D4", X"18", X"22", X"FE", X"FE", --3F90
  X"20", X"04", X"3E", X"D3", X"18", X"1A", X"FE", X"FD", --3F98
  X"20", X"04", X"3E", X"CE", X"18", X"12", X"FE", X"FC", --3FA0
  X"20", X"04", X"3E", X"ED", X"18", X"0A", X"FE", X"FB", --3FA8
  X"20", X"04", X"3E", X"EC", X"18", X"02", X"D6", X"56", --3FB0
  X"37", X"C9", X"46", X"23", X"7E", X"12", X"13", X"23", --3FB8
  X"10", X"FA", X"C9", X"FE", X"30", X"3F", X"D0", X"FE", --3FC0
  X"3A", X"D0", X"D6", X"30", X"37", X"C9", X"C5", X"D5", --3FC8
  X"46", X"23", X"BE", X"23", X"5E", X"23", X"56", X"28", --3FD0
  X"08", X"23", X"10", X"F6", X"37", X"3F", X"D1", X"C1", --3FD8
  X"C9", X"EB", X"D1", X"C1", X"CD", X"EE", X"3F", X"38", --3FE0
  X"02", X"BF", X"C9", X"BF", X"37", X"C9", X"E9", X"00", --3FE8
  X"4D", X"42", X"00", X"53", X"42", X"00", X"41", X"43", --3FF0
  X"00", X"52", X"47", X"00", X"4B", X"4D", X"00", X"01", --3FF8
  X"F3", X"01", X"00", X"40", X"61", X"C3", X"E1", X"3B", --4000
  X"2A", X"5D", X"5C", X"22", X"5F", X"5C", X"18", X"43", --4008
  X"C3", X"F2", X"15", X"FF", X"FF", X"FF", X"FF", X"FF", --4010
  X"2A", X"5D", X"5C", X"7E", X"CD", X"7D", X"00", X"D0", --4018
  X"CD", X"74", X"00", X"18", X"F7", X"FF", X"FF", X"FF", --4020
  X"C3", X"5B", X"33", X"FF", X"FF", X"FF", X"FF", X"FF", --4028
  X"C5", X"2A", X"61", X"5C", X"E5", X"C3", X"9E", X"16", --4030
  X"F5", X"E5", X"2A", X"78", X"5C", X"23", X"22", X"78", --4038
  X"5C", X"7C", X"B5", X"20", X"03", X"FD", X"34", X"40", --4040
  X"C5", X"D5", X"CD", X"6E", X"38", X"D1", X"C1", X"E1", --4048
  X"F1", X"FB", X"C9", X"E1", X"6E", X"FD", X"75", X"00", --4050
  X"ED", X"7B", X"3D", X"5C", X"C3", X"C5", X"16", X"FF", --4058
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F5", X"E5", --4060
  X"2A", X"B0", X"5C", X"7C", X"B5", X"20", X"01", X"E9", --4068
  X"E1", X"F1", X"ED", X"45", X"2A", X"5D", X"5C", X"23", --4070
  X"22", X"5D", X"5C", X"7E", X"C9", X"FE", X"21", X"D0", --4078
  X"FE", X"0D", X"C8", X"FE", X"10", X"D8", X"FE", X"18", --4080
  X"3F", X"D8", X"23", X"FE", X"16", X"38", X"01", X"23", --4088
  X"37", X"22", X"5D", X"5C", X"C9", X"BF", X"52", X"4E", --4090
  X"C4", X"49", X"4E", X"4B", X"45", X"59", X"A4", X"50", --4098
  X"C9", X"46", X"CE", X"50", X"4F", X"49", X"4E", X"D4", --40A0
  X"53", X"43", X"52", X"45", X"45", X"4E", X"A4", X"41", --40A8
  X"54", X"54", X"D2", X"41", X"D4", X"54", X"41", X"C2", --40B0
  X"56", X"41", X"4C", X"A4", X"43", X"4F", X"44", X"C5", --40B8
  X"56", X"41", X"CC", X"4C", X"45", X"CE", X"53", X"49", --40C0
  X"CE", X"43", X"4F", X"D3", X"54", X"41", X"CE", X"41", --40C8
  X"53", X"CE", X"41", X"43", X"D3", X"41", X"54", X"CE", --40D0
  X"4C", X"CE", X"45", X"58", X"D0", X"49", X"4E", X"D4", --40D8
  X"53", X"51", X"D2", X"53", X"47", X"CE", X"41", X"42", --40E0
  X"D3", X"50", X"45", X"45", X"CB", X"49", X"CE", X"55", --40E8
  X"53", X"D2", X"53", X"54", X"52", X"A4", X"43", X"48", --40F0
  X"52", X"A4", X"4E", X"4F", X"D4", X"42", X"49", X"CE", --40F8
  X"4F", X"D2", X"41", X"4E", X"C4", X"3C", X"BD", X"3E", --4100
  X"BD", X"3C", X"BE", X"4C", X"49", X"4E", X"C5", X"54", --4108
  X"48", X"45", X"CE", X"54", X"CF", X"53", X"54", X"45", --4110
  X"D0", X"44", X"45", X"46", X"20", X"46", X"CE", X"43", --4118
  X"41", X"D4", X"46", X"4F", X"52", X"4D", X"41", X"D4", --4120
  X"4D", X"4F", X"56", X"C5", X"45", X"52", X"41", X"53", --4128
  X"C5", X"4F", X"50", X"45", X"4E", X"20", X"A3", X"43", --4130
  X"4C", X"4F", X"53", X"45", X"20", X"A3", X"4D", X"45", --4138
  X"52", X"47", X"C5", X"56", X"45", X"52", X"49", X"46", --4140
  X"D9", X"42", X"45", X"45", X"D0", X"43", X"49", X"52", --4148
  X"43", X"4C", X"C5", X"49", X"4E", X"CB", X"50", X"41", --4150
  X"50", X"45", X"D2", X"46", X"4C", X"41", X"53", X"C8", --4158
  X"42", X"52", X"49", X"47", X"48", X"D4", X"49", X"4E", --4160
  X"56", X"45", X"52", X"53", X"C5", X"4F", X"56", X"45", --4168
  X"D2", X"4F", X"55", X"D4", X"4C", X"50", X"52", X"49", --4170
  X"4E", X"D4", X"4C", X"4C", X"49", X"53", X"D4", X"53", --4178
  X"54", X"4F", X"D0", X"52", X"45", X"41", X"C4", X"44", --4180
  X"41", X"54", X"C1", X"52", X"45", X"53", X"54", X"4F", --4188
  X"52", X"C5", X"4E", X"45", X"D7", X"42", X"4F", X"52", --4190
  X"44", X"45", X"D2", X"43", X"4F", X"4E", X"54", X"49", --4198
  X"4E", X"55", X"C5", X"44", X"49", X"CD", X"52", X"45", --41A0
  X"CD", X"46", X"4F", X"D2", X"47", X"4F", X"20", X"54", --41A8
  X"CF", X"47", X"4F", X"20", X"53", X"55", X"C2", X"49", --41B0
  X"4E", X"50", X"55", X"D4", X"4C", X"4F", X"41", X"C4", --41B8
  X"4C", X"49", X"53", X"D4", X"4C", X"45", X"D4", X"50", --41C0
  X"41", X"55", X"53", X"C5", X"4E", X"45", X"58", X"D4", --41C8
  X"50", X"4F", X"4B", X"C5", X"50", X"52", X"49", X"4E", --41D0
  X"D4", X"50", X"4C", X"4F", X"D4", X"52", X"55", X"CE", --41D8
  X"53", X"41", X"56", X"C5", X"52", X"41", X"4E", X"44", --41E0
  X"4F", X"4D", X"49", X"5A", X"C5", X"49", X"C6", X"43", --41E8
  X"4C", X"D3", X"44", X"52", X"41", X"D7", X"43", X"4C", --41F0
  X"45", X"41", X"D2", X"52", X"45", X"54", X"55", X"52", --41F8
  X"CE", X"43", X"4F", X"50", X"D9", X"42", X"48", X"59", --4200
  X"36", X"35", X"54", X"47", X"56", X"4E", X"4A", X"55", --4208
  X"37", X"34", X"52", X"46", X"43", X"4D", X"4B", X"49", --4210
  X"38", X"33", X"45", X"44", X"58", X"0E", X"4C", X"4F", --4218
  X"39", X"32", X"57", X"53", X"5A", X"20", X"0D", X"50", --4220
  X"30", X"31", X"51", X"41", X"E3", X"C4", X"E0", X"E4", --4228
  X"B4", X"BC", X"BD", X"BB", X"AF", X"B0", X"B1", X"C0", --4230
  X"A7", X"A6", X"BE", X"AD", X"B2", X"BA", X"E5", X"A5", --4238
  X"C2", X"E1", X"B3", X"B9", X"C1", X"B8", X"7E", X"DC", --4240
  X"DA", X"5C", X"B7", X"7B", X"7D", X"D8", X"BF", X"AE", --4248
  X"AA", X"AB", X"DD", X"DE", X"DF", X"7F", X"B5", X"D6", --4250
  X"7C", X"D5", X"5D", X"DB", X"B6", X"D9", X"5B", X"D7", --4258
  X"0C", X"07", X"06", X"04", X"05", X"08", X"0A", X"0B", --4260
  X"09", X"0F", X"E2", X"2A", X"3F", X"CD", X"C8", X"CC", --4268
  X"CB", X"5E", X"AC", X"2D", X"2B", X"3D", X"2E", X"2C", --4270
  X"3B", X"22", X"C7", X"3C", X"C3", X"3E", X"C5", X"2F", --4278
  X"C9", X"60", X"C6", X"3A", X"D0", X"CE", X"A8", X"CA", --4280
  X"D3", X"D4", X"D1", X"D2", X"A9", X"CF", X"2E", X"2F", --4288
  X"11", X"FF", X"FF", X"01", X"FE", X"FE", X"ED", X"78", --4290
  X"2F", X"E6", X"1F", X"28", X"0E", X"67", X"7D", X"14", --4298
  X"C0", X"D6", X"08", X"CB", X"3C", X"30", X"FA", X"53", --42A0
  X"5F", X"20", X"F4", X"2D", X"CB", X"00", X"38", X"E6", --42A8
  X"7A", X"3C", X"C8", X"FE", X"28", X"C8", X"FE", X"19", --42B0
  X"C8", X"7B", X"5A", X"57", X"FE", X"18", X"C9", X"CD", --42B8
  X"8E", X"02", X"C0", X"21", X"00", X"5C", X"CB", X"7E", --42C0
  X"20", X"07", X"23", X"35", X"2B", X"20", X"02", X"36", --42C8
  X"FF", X"7D", X"21", X"04", X"5C", X"BD", X"20", X"EE", --42D0
  X"CD", X"1E", X"03", X"D0", X"21", X"00", X"5C", X"BE", --42D8
  X"28", X"2E", X"EB", X"21", X"04", X"5C", X"BE", X"28", --42E0
  X"27", X"CB", X"7E", X"20", X"04", X"EB", X"CB", X"7E", --42E8
  X"C8", X"5F", X"77", X"23", X"36", X"05", X"23", X"3A", --42F0
  X"09", X"5C", X"77", X"23", X"FD", X"4E", X"07", X"FD", --42F8
  X"56", X"01", X"E5", X"CD", X"33", X"03", X"E1", X"77", --4300
  X"32", X"08", X"5C", X"FD", X"CB", X"01", X"EE", X"C9", --4308
  X"23", X"36", X"05", X"23", X"35", X"C0", X"3A", X"0A", --4310
  X"5C", X"77", X"23", X"7E", X"18", X"EA", X"42", X"16", --4318
  X"00", X"7B", X"FE", X"27", X"D0", X"FE", X"18", X"20", --4320
  X"03", X"CB", X"78", X"C0", X"21", X"05", X"02", X"19", --4328
  X"7E", X"37", X"C9", X"7B", X"FE", X"3A", X"38", X"2F", --4330
  X"0D", X"FA", X"4F", X"03", X"28", X"03", X"C6", X"4F", --4338
  X"C9", X"21", X"EB", X"01", X"04", X"28", X"03", X"21", --4340
  X"05", X"02", X"16", X"00", X"19", X"7E", X"C9", X"21", --4348
  X"29", X"02", X"CB", X"40", X"28", X"F4", X"CB", X"5A", --4350
  X"28", X"0A", X"FD", X"CB", X"30", X"5E", X"C0", X"04", --4358
  X"C0", X"C6", X"20", X"C9", X"C6", X"A5", X"C9", X"FE", --4360
  X"30", X"D8", X"0D", X"FA", X"9D", X"03", X"20", X"19", --4368
  X"21", X"54", X"02", X"CB", X"68", X"28", X"D3", X"FE", --4370
  X"38", X"30", X"07", X"D6", X"20", X"04", X"C8", X"C6", --4378
  X"08", X"C9", X"D6", X"36", X"04", X"C8", X"C6", X"FE", --4380
  X"C9", X"21", X"30", X"02", X"FE", X"39", X"28", X"BA", --4388
  X"FE", X"30", X"28", X"B6", X"E6", X"07", X"C6", X"80", --4390
  X"04", X"C8", X"EE", X"0F", X"C9", X"04", X"C8", X"CB", --4398
  X"68", X"21", X"30", X"02", X"20", X"A4", X"D6", X"10", --43A0
  X"FE", X"22", X"28", X"06", X"FE", X"20", X"C0", X"3E", --43A8
  X"5F", X"C9", X"3E", X"40", X"C9", X"F3", X"7D", X"CB", --43B0
  X"3D", X"CB", X"3D", X"2F", X"E6", X"03", X"4F", X"06", --43B8
  X"00", X"DD", X"21", X"D1", X"03", X"DD", X"09", X"3A", --43C0
  X"48", X"5C", X"E6", X"38", X"0F", X"0F", X"0F", X"F6", --43C8
  X"08", X"00", X"00", X"00", X"04", X"0C", X"0D", X"20", --43D0
  X"FD", X"0E", X"3F", X"05", X"C2", X"D6", X"03", X"EE", --43D8
  X"10", X"D3", X"FE", X"44", X"4F", X"CB", X"67", X"20", --43E0
  X"09", X"7A", X"B3", X"28", X"09", X"79", X"4D", X"1B", --43E8
  X"DD", X"E9", X"4D", X"0C", X"DD", X"E9", X"FB", X"C9", --43F0
  X"EF", X"31", X"27", X"C0", X"03", X"34", X"EC", X"6C", --43F8
  X"98", X"1F", X"F5", X"04", X"A1", X"0F", X"38", X"21", --4400
  X"92", X"5C", X"7E", X"A7", X"20", X"5E", X"23", X"4E", --4408
  X"23", X"46", X"78", X"17", X"9F", X"B9", X"20", X"54", --4410
  X"23", X"BE", X"20", X"50", X"78", X"C6", X"3C", X"F2", --4418
  X"25", X"04", X"E2", X"6C", X"04", X"06", X"FA", X"04", --4420
  X"D6", X"0C", X"30", X"FB", X"C6", X"0C", X"C5", X"21", --4428
  X"6E", X"04", X"CD", X"06", X"34", X"CD", X"B4", X"33", --4430
  X"EF", X"04", X"38", X"F1", X"86", X"77", X"EF", X"C0", --4438
  X"02", X"31", X"38", X"CD", X"94", X"1E", X"FE", X"0B", --4440
  X"30", X"22", X"EF", X"E0", X"04", X"E0", X"34", X"80", --4448
  X"43", X"55", X"9F", X"80", X"01", X"05", X"34", X"35", --4450
  X"71", X"03", X"38", X"CD", X"99", X"1E", X"C5", X"CD", --4458
  X"99", X"1E", X"E1", X"50", X"59", X"7A", X"B3", X"C8", --4460
  X"1B", X"C3", X"B5", X"03", X"CF", X"0A", X"89", X"02", --4468
  X"D0", X"12", X"86", X"89", X"0A", X"97", X"60", X"75", --4470
  X"89", X"12", X"D5", X"17", X"1F", X"89", X"1B", X"90", --4478
  X"41", X"02", X"89", X"24", X"D0", X"53", X"CA", X"89", --4480
  X"2E", X"9D", X"36", X"B1", X"89", X"38", X"FF", X"49", --4488
  X"3E", X"89", X"43", X"FF", X"6A", X"73", X"89", X"4F", --4490
  X"A7", X"00", X"54", X"89", X"5C", X"00", X"00", X"00", --4498
  X"89", X"69", X"14", X"F6", X"24", X"89", X"76", X"F1", --44A0
  X"10", X"05", X"CD", X"FB", X"24", X"3A", X"3B", X"5C", --44A8
  X"87", X"FA", X"8A", X"1C", X"E1", X"D0", X"E5", X"CD", --44B0
  X"F1", X"2B", X"62", X"6B", X"0D", X"F8", X"09", X"CB", --44B8
  X"FE", X"C9", X"21", X"3F", X"05", X"E5", X"21", X"80", --44C0
  X"1F", X"CB", X"7F", X"28", X"03", X"21", X"98", X"0C", --44C8
  X"08", X"13", X"DD", X"2B", X"F3", X"3E", X"02", X"47", --44D0
  X"10", X"FE", X"D3", X"FE", X"EE", X"0F", X"06", X"A4", --44D8
  X"2D", X"20", X"F5", X"05", X"25", X"F2", X"D8", X"04", --44E0
  X"06", X"2F", X"10", X"FE", X"D3", X"FE", X"3E", X"0D", --44E8
  X"06", X"37", X"10", X"FE", X"D3", X"FE", X"01", X"0E", --44F0
  X"3B", X"08", X"6F", X"C3", X"07", X"05", X"7A", X"B3", --44F8
  X"28", X"0C", X"DD", X"6E", X"00", X"7C", X"AD", X"67", --4500
  X"3E", X"01", X"37", X"C3", X"25", X"05", X"6C", X"18", --4508
  X"F4", X"79", X"CB", X"78", X"10", X"FE", X"30", X"04", --4510
  X"06", X"42", X"10", X"FE", X"D3", X"FE", X"06", X"3E", --4518
  X"20", X"EF", X"05", X"AF", X"3C", X"CB", X"15", X"C2", --4520
  X"14", X"05", X"1B", X"DD", X"23", X"06", X"31", X"3E", --4528
  X"7F", X"DB", X"FE", X"1F", X"D0", X"7A", X"3C", X"C2", --4530
  X"FE", X"04", X"06", X"3B", X"10", X"FE", X"C9", X"F5", --4538
  X"3A", X"48", X"5C", X"E6", X"38", X"0F", X"0F", X"0F", --4540
  X"D3", X"FE", X"3E", X"7F", X"DB", X"FE", X"1F", X"FB", --4548
  X"38", X"02", X"CF", X"0C", X"F1", X"C9", X"14", X"08", --4550
  X"15", X"F3", X"3E", X"0F", X"D3", X"FE", X"21", X"3F", --4558
  X"05", X"E5", X"DB", X"FE", X"1F", X"E6", X"20", X"F6", --4560
  X"02", X"4F", X"BF", X"C0", X"CD", X"E7", X"05", X"30", --4568
  X"FA", X"21", X"15", X"04", X"10", X"FE", X"2B", X"7C", --4570
  X"B5", X"20", X"F9", X"CD", X"E3", X"05", X"30", X"EB", --4578
  X"06", X"9C", X"CD", X"E3", X"05", X"30", X"E4", X"3E", --4580
  X"C6", X"B8", X"30", X"E0", X"24", X"20", X"F1", X"06", --4588
  X"C9", X"CD", X"E7", X"05", X"30", X"D5", X"78", X"FE", --4590
  X"D4", X"30", X"F4", X"CD", X"E7", X"05", X"D0", X"79", --4598
  X"EE", X"03", X"4F", X"26", X"00", X"06", X"B0", X"18", --45A0
  X"1F", X"08", X"20", X"07", X"30", X"0F", X"DD", X"75", --45A8
  X"00", X"18", X"0F", X"CB", X"11", X"AD", X"C0", X"79", --45B0
  X"1F", X"4F", X"13", X"18", X"07", X"DD", X"7E", X"00", --45B8
  X"AD", X"C0", X"DD", X"23", X"1B", X"08", X"06", X"B2", --45C0
  X"2E", X"01", X"CD", X"E3", X"05", X"D0", X"3E", X"CB", --45C8
  X"B8", X"CB", X"15", X"06", X"B0", X"D2", X"CA", X"05", --45D0
  X"7C", X"AD", X"67", X"7A", X"B3", X"20", X"CA", X"7C", --45D8
  X"FE", X"01", X"C9", X"CD", X"E7", X"05", X"D0", X"3E", --45E0
  X"16", X"3D", X"20", X"FD", X"A7", X"04", X"C8", X"3E", --45E8
  X"7F", X"DB", X"FE", X"1F", X"D0", X"A9", X"E6", X"20", --45F0
  X"28", X"F3", X"79", X"2F", X"4F", X"E6", X"07", X"F6", --45F8
  X"08", X"D3", X"FE", X"37", X"C9", X"F1", X"3A", X"74", --4600
  X"5C", X"D6", X"E0", X"32", X"74", X"5C", X"CD", X"8C", --4608
  X"1C", X"CD", X"30", X"25", X"28", X"3C", X"01", X"11", --4610
  X"00", X"3A", X"74", X"5C", X"A7", X"28", X"02", X"0E", --4618
  X"22", X"F7", X"D5", X"DD", X"E1", X"06", X"0B", X"3E", --4620
  X"20", X"12", X"13", X"10", X"FC", X"DD", X"36", X"01", --4628
  X"FF", X"CD", X"F1", X"2B", X"21", X"F6", X"FF", X"0B", --4630
  X"09", X"03", X"30", X"0F", X"3A", X"74", X"5C", X"A7", --4638
  X"20", X"02", X"CF", X"0E", X"78", X"B1", X"28", X"0A", --4640
  X"01", X"0A", X"00", X"DD", X"E5", X"E1", X"23", X"EB", --4648
  X"ED", X"B0", X"DF", X"FE", X"E4", X"20", X"49", X"3A", --4650
  X"74", X"5C", X"FE", X"03", X"CA", X"8A", X"1C", X"E7", --4658
  X"CD", X"B2", X"28", X"CB", X"F9", X"30", X"0B", X"21", --4660
  X"00", X"00", X"3A", X"74", X"5C", X"3D", X"28", X"15", --4668
  X"CF", X"01", X"C2", X"8A", X"1C", X"CD", X"30", X"25", --4670
  X"28", X"18", X"23", X"7E", X"DD", X"77", X"0B", X"23", --4678
  X"7E", X"DD", X"77", X"0C", X"23", X"DD", X"71", X"0E", --4680
  X"3E", X"01", X"CB", X"71", X"28", X"01", X"3C", X"DD", --4688
  X"77", X"00", X"EB", X"E7", X"FE", X"29", X"20", X"DA", --4690
  X"E7", X"CD", X"EE", X"1B", X"EB", X"C3", X"5A", X"07", --4698
  X"FE", X"AA", X"20", X"1F", X"3A", X"74", X"5C", X"FE", --46A0
  X"03", X"CA", X"8A", X"1C", X"E7", X"CD", X"EE", X"1B", --46A8
  X"DD", X"36", X"0B", X"00", X"DD", X"36", X"0C", X"1B", --46B0
  X"21", X"00", X"40", X"DD", X"75", X"0D", X"DD", X"74", --46B8
  X"0E", X"18", X"4D", X"FE", X"AF", X"20", X"4F", X"3A", --46C0
  X"74", X"5C", X"FE", X"03", X"CA", X"8A", X"1C", X"E7", --46C8
  X"CD", X"48", X"20", X"20", X"0C", X"3A", X"74", X"5C", --46D0
  X"A7", X"CA", X"8A", X"1C", X"CD", X"E6", X"1C", X"18", --46D8
  X"0F", X"CD", X"82", X"1C", X"DF", X"FE", X"2C", X"28", --46E0
  X"0C", X"3A", X"74", X"5C", X"A7", X"CA", X"8A", X"1C", --46E8
  X"CD", X"E6", X"1C", X"18", X"04", X"E7", X"CD", X"82", --46F0
  X"1C", X"CD", X"EE", X"1B", X"CD", X"99", X"1E", X"DD", --46F8
  X"71", X"0B", X"DD", X"70", X"0C", X"CD", X"99", X"1E", --4700
  X"DD", X"71", X"0D", X"DD", X"70", X"0E", X"60", X"69", --4708
  X"DD", X"36", X"00", X"03", X"18", X"44", X"FE", X"CA", --4710
  X"28", X"09", X"CD", X"EE", X"1B", X"DD", X"36", X"0E", --4718
  X"80", X"18", X"17", X"3A", X"74", X"5C", X"A7", X"C2", --4720
  X"8A", X"1C", X"E7", X"CD", X"82", X"1C", X"CD", X"EE", --4728
  X"1B", X"CD", X"99", X"1E", X"DD", X"71", X"0D", X"DD", --4730
  X"70", X"0E", X"DD", X"36", X"00", X"00", X"2A", X"59", --4738
  X"5C", X"ED", X"5B", X"53", X"5C", X"37", X"ED", X"52", --4740
  X"DD", X"75", X"0B", X"DD", X"74", X"0C", X"2A", X"4B", --4748
  X"5C", X"ED", X"52", X"DD", X"75", X"0F", X"DD", X"74", --4750
  X"10", X"EB", X"3A", X"74", X"5C", X"A7", X"CA", X"70", --4758
  X"09", X"E5", X"01", X"11", X"00", X"DD", X"09", X"DD", --4760
  X"E5", X"11", X"11", X"00", X"AF", X"37", X"CD", X"56", --4768
  X"05", X"DD", X"E1", X"30", X"F2", X"3E", X"FE", X"CD", --4770
  X"01", X"16", X"FD", X"36", X"52", X"03", X"0E", X"80", --4778
  X"DD", X"7E", X"00", X"DD", X"BE", X"EF", X"20", X"02", --4780
  X"0E", X"F6", X"FE", X"04", X"30", X"D9", X"11", X"C0", --4788
  X"09", X"C5", X"CD", X"0A", X"0C", X"C1", X"DD", X"E5", --4790
  X"D1", X"21", X"F0", X"FF", X"19", X"06", X"0A", X"7E", --4798
  X"3C", X"20", X"03", X"79", X"80", X"4F", X"13", X"1A", --47A0
  X"BE", X"23", X"20", X"01", X"0C", X"D7", X"10", X"F6", --47A8
  X"CB", X"79", X"20", X"B3", X"3E", X"0D", X"D7", X"E1", --47B0
  X"DD", X"7E", X"00", X"FE", X"03", X"28", X"0C", X"3A", --47B8
  X"74", X"5C", X"3D", X"CA", X"08", X"08", X"FE", X"02", --47C0
  X"CA", X"B6", X"08", X"E5", X"DD", X"6E", X"FA", X"DD", --47C8
  X"66", X"FB", X"DD", X"5E", X"0B", X"DD", X"56", X"0C", --47D0
  X"7C", X"B5", X"28", X"0D", X"ED", X"52", X"38", X"26", --47D8
  X"28", X"07", X"DD", X"7E", X"00", X"FE", X"03", X"20", --47E0
  X"1D", X"E1", X"7C", X"B5", X"20", X"06", X"DD", X"6E", --47E8
  X"0D", X"DD", X"66", X"0E", X"E5", X"DD", X"E1", X"3A", --47F0
  X"74", X"5C", X"FE", X"02", X"37", X"20", X"01", X"A7", --47F8
  X"3E", X"FF", X"CD", X"56", X"05", X"D8", X"CF", X"1A", --4800
  X"DD", X"5E", X"0B", X"DD", X"56", X"0C", X"E5", X"7C", --4808
  X"B5", X"20", X"06", X"13", X"13", X"13", X"EB", X"18", --4810
  X"0C", X"DD", X"6E", X"FA", X"DD", X"66", X"FB", X"EB", --4818
  X"37", X"ED", X"52", X"38", X"09", X"11", X"05", X"00", --4820
  X"19", X"44", X"4D", X"CD", X"05", X"1F", X"E1", X"DD", --4828
  X"7E", X"00", X"A7", X"28", X"3E", X"7C", X"B5", X"28", --4830
  X"13", X"2B", X"46", X"2B", X"4E", X"2B", X"03", X"03", --4838
  X"03", X"DD", X"22", X"5F", X"5C", X"CD", X"E8", X"19", --4840
  X"DD", X"2A", X"5F", X"5C", X"2A", X"59", X"5C", X"2B", --4848
  X"DD", X"4E", X"0B", X"DD", X"46", X"0C", X"C5", X"03", --4850
  X"03", X"03", X"DD", X"7E", X"FD", X"F5", X"CD", X"55", --4858
  X"16", X"23", X"F1", X"77", X"D1", X"23", X"73", X"23", --4860
  X"72", X"23", X"E5", X"DD", X"E1", X"37", X"3E", X"FF", --4868
  X"C3", X"02", X"08", X"EB", X"2A", X"59", X"5C", X"2B", --4870
  X"DD", X"22", X"5F", X"5C", X"DD", X"4E", X"0B", X"DD", --4878
  X"46", X"0C", X"C5", X"CD", X"E5", X"19", X"C1", X"E5", --4880
  X"C5", X"CD", X"55", X"16", X"DD", X"2A", X"5F", X"5C", --4888
  X"23", X"DD", X"4E", X"0F", X"DD", X"46", X"10", X"09", --4890
  X"22", X"4B", X"5C", X"DD", X"66", X"0E", X"7C", X"E6", --4898
  X"C0", X"20", X"0A", X"DD", X"6E", X"0D", X"22", X"42", --48A0
  X"5C", X"FD", X"36", X"0A", X"00", X"D1", X"DD", X"E1", --48A8
  X"37", X"3E", X"FF", X"C3", X"02", X"08", X"DD", X"4E", --48B0
  X"0B", X"DD", X"46", X"0C", X"C5", X"03", X"F7", X"36", --48B8
  X"80", X"EB", X"D1", X"E5", X"E5", X"DD", X"E1", X"37", --48C0
  X"3E", X"FF", X"CD", X"02", X"08", X"E1", X"ED", X"5B", --48C8
  X"53", X"5C", X"7E", X"E6", X"C0", X"20", X"19", X"1A", --48D0
  X"13", X"BE", X"23", X"20", X"02", X"1A", X"BE", X"1B", --48D8
  X"2B", X"30", X"08", X"E5", X"EB", X"CD", X"B8", X"19", --48E0
  X"E1", X"18", X"EC", X"CD", X"2C", X"09", X"18", X"E2", --48E8
  X"7E", X"4F", X"FE", X"80", X"C8", X"E5", X"2A", X"4B", --48F0
  X"5C", X"7E", X"FE", X"80", X"28", X"25", X"B9", X"28", --48F8
  X"08", X"C5", X"CD", X"B8", X"19", X"C1", X"EB", X"18", --4900
  X"F0", X"E6", X"E0", X"FE", X"A0", X"20", X"12", X"D1", --4908
  X"D5", X"E5", X"23", X"13", X"1A", X"BE", X"20", X"06", --4910
  X"17", X"30", X"F7", X"E1", X"18", X"03", X"E1", X"18", --4918
  X"E0", X"3E", X"FF", X"D1", X"EB", X"3C", X"37", X"CD", --4920
  X"2C", X"09", X"18", X"C4", X"20", X"10", X"08", X"22", --4928
  X"5F", X"5C", X"EB", X"CD", X"B8", X"19", X"CD", X"E8", --4930
  X"19", X"EB", X"2A", X"5F", X"5C", X"08", X"08", X"D5", --4938
  X"CD", X"B8", X"19", X"22", X"5F", X"5C", X"2A", X"53", --4940
  X"5C", X"E3", X"C5", X"08", X"38", X"07", X"2B", X"CD", --4948
  X"55", X"16", X"23", X"18", X"03", X"CD", X"55", X"16", --4950
  X"23", X"C1", X"D1", X"ED", X"53", X"53", X"5C", X"ED", --4958
  X"5B", X"5F", X"5C", X"C5", X"D5", X"EB", X"ED", X"B0", --4960
  X"E1", X"C1", X"D5", X"CD", X"E8", X"19", X"D1", X"C9", --4968
  X"E5", X"3E", X"FD", X"CD", X"01", X"16", X"AF", X"11", --4970
  X"A1", X"09", X"CD", X"0A", X"0C", X"FD", X"CB", X"02", --4978
  X"EE", X"CD", X"D4", X"15", X"DD", X"E5", X"11", X"11", --4980
  X"00", X"AF", X"CD", X"C2", X"04", X"DD", X"E1", X"06", --4988
  X"32", X"76", X"10", X"FD", X"DD", X"5E", X"0B", X"DD", --4990
  X"56", X"0C", X"3E", X"FF", X"DD", X"E1", X"C3", X"C2", --4998
  X"04", X"80", X"53", X"74", X"61", X"72", X"74", X"20", --49A0
  X"74", X"61", X"70", X"65", X"2C", X"20", X"74", X"68", --49A8
  X"65", X"6E", X"20", X"70", X"72", X"65", X"73", X"73", --49B0
  X"20", X"61", X"6E", X"79", X"20", X"6B", X"65", X"79", --49B8
  X"AE", X"0D", X"50", X"72", X"6F", X"67", X"72", X"61", --49C0
  X"6D", X"3A", X"A0", X"0D", X"4E", X"75", X"6D", X"62", --49C8
  X"65", X"72", X"20", X"61", X"72", X"72", X"61", X"79", --49D0
  X"3A", X"A0", X"0D", X"43", X"68", X"61", X"72", X"61", --49D8
  X"63", X"74", X"65", X"72", X"20", X"61", X"72", X"72", --49E0
  X"61", X"79", X"3A", X"A0", X"0D", X"42", X"79", X"74", --49E8
  X"65", X"73", X"3A", X"A0", X"CD", X"03", X"0B", X"FE", --49F0
  X"20", X"D2", X"D9", X"0A", X"FE", X"06", X"38", X"69", --49F8
  X"FE", X"18", X"30", X"65", X"21", X"0B", X"0A", X"5F", --4A00
  X"16", X"00", X"19", X"5E", X"19", X"E5", X"C3", X"03", --4A08
  X"0B", X"4E", X"57", X"10", X"29", X"54", X"53", X"52", --4A10
  X"37", X"50", X"4F", X"5F", X"5E", X"5D", X"5C", X"5B", --4A18
  X"5A", X"54", X"53", X"0C", X"3E", X"22", X"B9", X"20", --4A20
  X"11", X"FD", X"CB", X"01", X"4E", X"20", X"09", X"04", --4A28
  X"0E", X"02", X"3E", X"18", X"B8", X"20", X"03", X"05", --4A30
  X"0E", X"21", X"C3", X"D9", X"0D", X"3A", X"91", X"5C", --4A38
  X"F5", X"FD", X"36", X"57", X"01", X"3E", X"20", X"CD", --4A40
  X"65", X"0B", X"F1", X"32", X"91", X"5C", X"C9", X"FD", --4A48
  X"CB", X"01", X"4E", X"C2", X"CD", X"0E", X"0E", X"21", --4A50
  X"CD", X"55", X"0C", X"05", X"C3", X"D9", X"0D", X"CD", --4A58
  X"03", X"0B", X"79", X"3D", X"3D", X"E6", X"10", X"18", --4A60
  X"5A", X"3E", X"3F", X"18", X"6C", X"11", X"87", X"0A", --4A68
  X"32", X"0F", X"5C", X"18", X"0B", X"11", X"6D", X"0A", --4A70
  X"18", X"03", X"11", X"87", X"0A", X"32", X"0E", X"5C", --4A78
  X"2A", X"51", X"5C", X"73", X"23", X"72", X"C9", X"11", --4A80
  X"F4", X"09", X"CD", X"80", X"0A", X"2A", X"0E", X"5C", --4A88
  X"57", X"7D", X"FE", X"16", X"DA", X"11", X"22", X"20", --4A90
  X"29", X"44", X"4A", X"3E", X"1F", X"91", X"38", X"0C", --4A98
  X"C6", X"02", X"4F", X"FD", X"CB", X"01", X"4E", X"20", --4AA0
  X"16", X"3E", X"16", X"90", X"DA", X"9F", X"1E", X"3C", --4AA8
  X"47", X"04", X"FD", X"CB", X"02", X"46", X"C2", X"55", --4AB0
  X"0C", X"FD", X"BE", X"31", X"DA", X"86", X"0C", X"C3", --4AB8
  X"D9", X"0D", X"7C", X"CD", X"03", X"0B", X"81", X"3D", --4AC0
  X"E6", X"1F", X"C8", X"57", X"FD", X"CB", X"01", X"C6", --4AC8
  X"3E", X"20", X"CD", X"3B", X"0C", X"15", X"20", X"F8", --4AD0
  X"C9", X"CD", X"24", X"0B", X"FD", X"CB", X"01", X"4E", --4AD8
  X"20", X"1A", X"FD", X"CB", X"02", X"46", X"20", X"08", --4AE0
  X"ED", X"43", X"88", X"5C", X"22", X"84", X"5C", X"C9", --4AE8
  X"ED", X"43", X"8A", X"5C", X"ED", X"43", X"82", X"5C", --4AF0
  X"22", X"86", X"5C", X"C9", X"FD", X"71", X"45", X"22", --4AF8
  X"80", X"5C", X"C9", X"FD", X"CB", X"01", X"4E", X"20", --4B00
  X"14", X"ED", X"4B", X"88", X"5C", X"2A", X"84", X"5C", --4B08
  X"FD", X"CB", X"02", X"46", X"C8", X"ED", X"4B", X"8A", --4B10
  X"5C", X"2A", X"86", X"5C", X"C9", X"FD", X"4E", X"45", --4B18
  X"2A", X"80", X"5C", X"C9", X"FE", X"80", X"38", X"3D", --4B20
  X"FE", X"90", X"30", X"26", X"47", X"CD", X"38", X"0B", --4B28
  X"CD", X"03", X"0B", X"11", X"92", X"5C", X"18", X"47", --4B30
  X"21", X"92", X"5C", X"CD", X"3E", X"0B", X"CB", X"18", --4B38
  X"9F", X"E6", X"0F", X"4F", X"CB", X"18", X"9F", X"E6", --4B40
  X"F0", X"B1", X"0E", X"04", X"77", X"23", X"0D", X"20", --4B48
  X"FB", X"C9", X"C3", X"9F", X"3B", X"00", X"C6", X"15", --4B50
  X"C5", X"ED", X"4B", X"7B", X"5C", X"18", X"0B", X"CD", --4B58
  X"10", X"0C", X"C3", X"03", X"0B", X"C5", X"ED", X"4B", --4B60
  X"36", X"5C", X"EB", X"21", X"3B", X"5C", X"CB", X"86", --4B68
  X"FE", X"20", X"20", X"02", X"CB", X"C6", X"26", X"00", --4B70
  X"6F", X"29", X"29", X"29", X"09", X"C1", X"EB", X"79", --4B78
  X"3D", X"3E", X"21", X"20", X"0E", X"05", X"4F", X"FD", --4B80
  X"CB", X"01", X"4E", X"28", X"06", X"D5", X"CD", X"CD", --4B88
  X"0E", X"D1", X"79", X"B9", X"D5", X"CC", X"55", X"0C", --4B90
  X"D1", X"C5", X"E5", X"3A", X"91", X"5C", X"06", X"FF", --4B98
  X"1F", X"38", X"01", X"04", X"1F", X"1F", X"9F", X"4F", --4BA0
  X"3E", X"08", X"A7", X"FD", X"CB", X"01", X"4E", X"28", --4BA8
  X"05", X"FD", X"CB", X"30", X"CE", X"37", X"EB", X"08", --4BB0
  X"1A", X"A0", X"AE", X"A9", X"12", X"08", X"38", X"13", --4BB8
  X"14", X"23", X"3D", X"20", X"F2", X"EB", X"25", X"FD", --4BC0
  X"CB", X"01", X"4E", X"CC", X"DB", X"0B", X"E1", X"C1", --4BC8
  X"0D", X"23", X"C9", X"08", X"3E", X"20", X"83", X"5F", --4BD0
  X"08", X"18", X"E6", X"7C", X"0F", X"0F", X"0F", X"E6", --4BD8
  X"03", X"F6", X"58", X"67", X"ED", X"5B", X"8F", X"5C", --4BE0
  X"7E", X"AB", X"A2", X"AB", X"FD", X"CB", X"57", X"76", --4BE8
  X"28", X"08", X"E6", X"C7", X"CB", X"57", X"20", X"02", --4BF0
  X"EE", X"38", X"FD", X"CB", X"57", X"66", X"28", X"08", --4BF8
  X"E6", X"F8", X"CB", X"6F", X"20", X"02", X"EE", X"07", --4C00
  X"77", X"C9", X"E5", X"26", X"00", X"E3", X"18", X"04", --4C08
  X"11", X"95", X"00", X"F5", X"CD", X"41", X"0C", X"38", --4C10
  X"09", X"3E", X"20", X"FD", X"CB", X"01", X"46", X"CC", --4C18
  X"3B", X"0C", X"1A", X"E6", X"7F", X"CD", X"3B", X"0C", --4C20
  X"1A", X"13", X"87", X"30", X"F5", X"D1", X"FE", X"48", --4C28
  X"28", X"03", X"FE", X"82", X"D8", X"7A", X"FE", X"03", --4C30
  X"D8", X"3E", X"20", X"D5", X"D9", X"D7", X"D9", X"D1", --4C38
  X"C9", X"F5", X"EB", X"3C", X"CB", X"7E", X"23", X"28", --4C40
  X"FB", X"3D", X"20", X"F8", X"EB", X"F1", X"FE", X"20", --4C48
  X"D8", X"1A", X"D6", X"41", X"C9", X"FD", X"CB", X"01", --4C50
  X"4E", X"C0", X"11", X"D9", X"0D", X"D5", X"78", X"FD", --4C58
  X"CB", X"02", X"46", X"C2", X"02", X"0D", X"FD", X"BE", --4C60
  X"31", X"38", X"1B", X"C0", X"FD", X"CB", X"02", X"66", --4C68
  X"28", X"16", X"FD", X"5E", X"2D", X"1D", X"28", X"5A", --4C70
  X"3E", X"00", X"CD", X"01", X"16", X"ED", X"7B", X"3F", --4C78
  X"5C", X"FD", X"CB", X"02", X"A6", X"C9", X"CF", X"04", --4C80
  X"FD", X"35", X"52", X"20", X"45", X"3E", X"18", X"90", --4C88
  X"32", X"8C", X"5C", X"2A", X"8F", X"5C", X"E5", X"3A", --4C90
  X"91", X"5C", X"F5", X"3E", X"FD", X"CD", X"01", X"16", --4C98
  X"AF", X"11", X"F8", X"0C", X"CD", X"0A", X"0C", X"FD", --4CA0
  X"CB", X"02", X"EE", X"21", X"3B", X"5C", X"CB", X"DE", --4CA8
  X"CB", X"AE", X"D9", X"CD", X"D4", X"15", X"D9", X"FE", --4CB0
  X"20", X"28", X"45", X"FE", X"E2", X"28", X"41", X"F6", --4CB8
  X"20", X"FE", X"6E", X"28", X"3B", X"3E", X"FE", X"CD", --4CC0
  X"01", X"16", X"F1", X"32", X"91", X"5C", X"E1", X"22", --4CC8
  X"8F", X"5C", X"CD", X"FE", X"0D", X"FD", X"46", X"31", --4CD0
  X"04", X"0E", X"21", X"C5", X"CD", X"9B", X"0E", X"7C", --4CD8
  X"0F", X"0F", X"0F", X"E6", X"03", X"F6", X"58", X"67", --4CE0
  X"11", X"E0", X"5A", X"1A", X"4E", X"06", X"20", X"EB", --4CE8
  X"12", X"71", X"13", X"23", X"10", X"FA", X"C1", X"C9", --4CF0
  X"80", X"73", X"63", X"72", X"6F", X"6C", X"6C", X"BF", --4CF8
  X"CF", X"0C", X"FE", X"02", X"38", X"80", X"FD", X"86", --4D00
  X"31", X"D6", X"19", X"D0", X"ED", X"44", X"C5", X"47", --4D08
  X"2A", X"8F", X"5C", X"E5", X"2A", X"91", X"5C", X"E5", --4D10
  X"CD", X"4D", X"0D", X"78", X"F5", X"21", X"6B", X"5C", --4D18
  X"46", X"78", X"3C", X"77", X"21", X"89", X"5C", X"BE", --4D20
  X"38", X"03", X"34", X"06", X"18", X"CD", X"00", X"0E", --4D28
  X"F1", X"3D", X"20", X"E8", X"E1", X"FD", X"75", X"57", --4D30
  X"E1", X"22", X"8F", X"5C", X"ED", X"4B", X"88", X"5C", --4D38
  X"FD", X"CB", X"02", X"86", X"CD", X"D9", X"0D", X"FD", --4D40
  X"CB", X"02", X"C6", X"C1", X"C9", X"AF", X"2A", X"8D", --4D48
  X"5C", X"FD", X"CB", X"02", X"46", X"28", X"04", X"67", --4D50
  X"FD", X"6E", X"0E", X"22", X"8F", X"5C", X"21", X"91", --4D58
  X"5C", X"20", X"02", X"7E", X"0F", X"AE", X"E6", X"55", --4D60
  X"AE", X"77", X"C9", X"CD", X"AF", X"0D", X"21", X"3C", --4D68
  X"5C", X"CB", X"AE", X"CB", X"C6", X"CD", X"4D", X"0D", --4D70
  X"FD", X"46", X"31", X"CD", X"44", X"0E", X"21", X"C0", --4D78
  X"5A", X"3A", X"8D", X"5C", X"05", X"18", X"07", X"0E", --4D80
  X"20", X"2B", X"77", X"0D", X"20", X"FB", X"10", X"F7", --4D88
  X"FD", X"36", X"31", X"02", X"3E", X"FD", X"CD", X"01", --4D90
  X"16", X"2A", X"51", X"5C", X"11", X"F4", X"09", X"A7", --4D98
  X"73", X"23", X"72", X"23", X"11", X"A8", X"10", X"3F", --4DA0
  X"38", X"F6", X"01", X"21", X"17", X"18", X"2A", X"21", --4DA8
  X"00", X"00", X"22", X"7D", X"5C", X"FD", X"CB", X"30", --4DB0
  X"86", X"CD", X"94", X"0D", X"3E", X"FE", X"CD", X"01", --4DB8
  X"16", X"CD", X"4D", X"0D", X"06", X"18", X"CD", X"44", --4DC0
  X"0E", X"2A", X"51", X"5C", X"11", X"F4", X"09", X"73", --4DC8
  X"23", X"72", X"FD", X"36", X"52", X"01", X"01", X"21", --4DD0
  X"18", X"21", X"00", X"5B", X"FD", X"CB", X"01", X"4E", --4DD8
  X"20", X"12", X"78", X"FD", X"CB", X"02", X"46", X"28", --4DE0
  X"05", X"FD", X"86", X"31", X"D6", X"18", X"C5", X"47", --4DE8
  X"CD", X"9B", X"0E", X"C1", X"3E", X"21", X"91", X"5F", --4DF0
  X"16", X"00", X"19", X"C3", X"DC", X"0A", X"06", X"17", --4DF8
  X"CD", X"9B", X"0E", X"0E", X"08", X"C5", X"E5", X"78", --4E00
  X"E6", X"07", X"78", X"20", X"0C", X"EB", X"21", X"E0", --4E08
  X"F8", X"19", X"EB", X"01", X"20", X"00", X"3D", X"ED", --4E10
  X"B0", X"EB", X"21", X"E0", X"FF", X"19", X"EB", X"47", --4E18
  X"E6", X"07", X"0F", X"0F", X"0F", X"4F", X"78", X"06", --4E20
  X"00", X"ED", X"B0", X"06", X"07", X"09", X"E6", X"F8", --4E28
  X"20", X"DB", X"E1", X"24", X"C1", X"0D", X"20", X"CD", --4E30
  X"CD", X"88", X"0E", X"21", X"E0", X"FF", X"19", X"EB", --4E38
  X"ED", X"B0", X"06", X"01", X"C5", X"CD", X"9B", X"0E", --4E40
  X"0E", X"08", X"C5", X"E5", X"78", X"E6", X"07", X"0F", --4E48
  X"0F", X"0F", X"4F", X"78", X"06", X"00", X"0D", X"54", --4E50
  X"5D", X"36", X"00", X"13", X"ED", X"B0", X"11", X"01", --4E58
  X"07", X"19", X"3D", X"E6", X"F8", X"47", X"20", X"E5", --4E60
  X"E1", X"24", X"C1", X"0D", X"20", X"DC", X"CD", X"88", --4E68
  X"0E", X"62", X"6B", X"13", X"3A", X"8D", X"5C", X"FD", --4E70
  X"CB", X"02", X"46", X"28", X"03", X"3A", X"48", X"5C", --4E78
  X"77", X"0B", X"ED", X"B0", X"C1", X"0E", X"21", X"C9", --4E80
  X"7C", X"0F", X"0F", X"0F", X"3D", X"F6", X"50", X"67", --4E88
  X"EB", X"61", X"68", X"29", X"29", X"29", X"29", X"29", --4E90
  X"44", X"4D", X"C9", X"3E", X"18", X"90", X"57", X"0F", --4E98
  X"0F", X"0F", X"E6", X"E0", X"6F", X"7A", X"E6", X"18", --4EA0
  X"F6", X"40", X"67", X"C9", X"F3", X"06", X"B0", X"21", --4EA8
  X"00", X"40", X"E5", X"C5", X"CD", X"F4", X"0E", X"C1", --4EB0
  X"E1", X"24", X"7C", X"E6", X"07", X"20", X"0A", X"7D", --4EB8
  X"C6", X"20", X"6F", X"3F", X"9F", X"E6", X"F8", X"84", --4EC0
  X"67", X"10", X"E7", X"18", X"0D", X"F3", X"21", X"00", --4EC8
  X"5B", X"06", X"08", X"C5", X"CD", X"F4", X"0E", X"C1", --4ED0
  X"10", X"F9", X"3E", X"04", X"D3", X"FB", X"FB", X"21", --4ED8
  X"00", X"5B", X"FD", X"75", X"46", X"AF", X"47", X"77", --4EE0
  X"23", X"10", X"FC", X"FD", X"CB", X"30", X"8E", X"0E", --4EE8
  X"21", X"C3", X"D9", X"0D", X"78", X"FE", X"03", X"9F", --4EF0
  X"E6", X"02", X"D3", X"FB", X"57", X"CD", X"54", X"1F", --4EF8
  X"38", X"0A", X"3E", X"04", X"D3", X"FB", X"FB", X"CD", --4F00
  X"DF", X"0E", X"CF", X"0C", X"DB", X"FB", X"87", X"F8", --4F08
  X"30", X"EB", X"0E", X"20", X"5E", X"23", X"06", X"08", --4F10
  X"CB", X"12", X"CB", X"13", X"CB", X"1A", X"DB", X"FB", --4F18
  X"1F", X"30", X"FB", X"7A", X"D3", X"FB", X"10", X"F0", --4F20
  X"0D", X"20", X"E9", X"C9", X"2A", X"3D", X"5C", X"E5", --4F28
  X"21", X"7F", X"10", X"E5", X"ED", X"73", X"3D", X"5C", --4F30
  X"CD", X"D4", X"15", X"F5", X"16", X"00", X"FD", X"5E", --4F38
  X"FF", X"21", X"C8", X"00", X"CD", X"B5", X"03", X"F1", --4F40
  X"21", X"38", X"0F", X"E5", X"FE", X"18", X"30", X"31", --4F48
  X"FE", X"07", X"38", X"2D", X"FE", X"10", X"38", X"3A", --4F50
  X"01", X"02", X"00", X"57", X"FE", X"16", X"38", X"0C", --4F58
  X"03", X"FD", X"CB", X"37", X"7E", X"CA", X"1E", X"10", --4F60
  X"CD", X"D4", X"15", X"5F", X"CD", X"D4", X"15", X"D5", --4F68
  X"2A", X"5B", X"5C", X"FD", X"CB", X"07", X"86", X"CD", --4F70
  X"55", X"16", X"C1", X"23", X"70", X"23", X"71", X"18", --4F78
  X"0A", X"FD", X"CB", X"07", X"86", X"2A", X"5B", X"5C", --4F80
  X"CD", X"52", X"16", X"12", X"13", X"ED", X"53", X"5B", --4F88
  X"5C", X"C9", X"5F", X"16", X"00", X"21", X"99", X"0F", --4F90
  X"19", X"5E", X"19", X"E5", X"2A", X"5B", X"5C", X"C9", --4F98
  X"09", X"66", X"6A", X"50", X"B5", X"70", X"7E", X"CF", --4FA0
  X"D4", X"2A", X"49", X"5C", X"FD", X"CB", X"37", X"6E", --4FA8
  X"C2", X"97", X"10", X"CD", X"6E", X"19", X"CD", X"95", --4FB0
  X"16", X"7A", X"B3", X"CA", X"97", X"10", X"E5", X"23", --4FB8
  X"4E", X"23", X"46", X"21", X"0A", X"00", X"09", X"44", --4FC0
  X"4D", X"CD", X"05", X"1F", X"CD", X"97", X"10", X"2A", --4FC8
  X"51", X"5C", X"E3", X"E5", X"3E", X"FF", X"CD", X"01", --4FD0
  X"16", X"E1", X"2B", X"FD", X"35", X"0F", X"CD", X"55", --4FD8
  X"18", X"FD", X"34", X"0F", X"2A", X"59", X"5C", X"23", --4FE0
  X"23", X"23", X"23", X"22", X"5B", X"5C", X"E1", X"CD", --4FE8
  X"15", X"16", X"C9", X"FD", X"CB", X"37", X"6E", X"20", --4FF0
  X"08", X"21", X"49", X"5C", X"CD", X"0F", X"19", X"18", --4FF8
  X"6D", X"FD", X"36", X"00", X"10", X"18", X"1D", X"CD", --5000
  X"31", X"10", X"18", X"05", X"7E", X"FE", X"0D", X"C8", --5008
  X"23", X"22", X"5B", X"5C", X"C9", X"CD", X"31", X"10", --5010
  X"01", X"01", X"00", X"C3", X"E8", X"19", X"CD", X"D4", --5018
  X"15", X"CD", X"D4", X"15", X"E1", X"E1", X"E1", X"22", --5020
  X"3D", X"5C", X"FD", X"CB", X"00", X"7E", X"C0", X"F9", --5028
  X"C9", X"37", X"CD", X"95", X"11", X"ED", X"52", X"19", --5030
  X"23", X"C1", X"D8", X"C5", X"44", X"4D", X"62", X"6B", --5038
  X"23", X"1A", X"E6", X"F0", X"FE", X"10", X"20", X"09", --5040
  X"23", X"1A", X"D6", X"17", X"CE", X"00", X"20", X"01", --5048
  X"23", X"A7", X"ED", X"42", X"09", X"EB", X"38", X"E6", --5050
  X"C9", X"FD", X"CB", X"37", X"6E", X"C0", X"2A", X"49", --5058
  X"5C", X"CD", X"6E", X"19", X"EB", X"CD", X"95", X"16", --5060
  X"21", X"4A", X"5C", X"CD", X"1C", X"19", X"CD", X"95", --5068
  X"17", X"3E", X"00", X"C3", X"01", X"16", X"FD", X"CB", --5070
  X"37", X"7E", X"28", X"A8", X"C3", X"81", X"0F", X"FD", --5078
  X"CB", X"30", X"66", X"28", X"A1", X"FD", X"36", X"00", --5080
  X"FF", X"16", X"00", X"FD", X"5E", X"FE", X"21", X"90", --5088
  X"1A", X"CD", X"B5", X"03", X"C3", X"30", X"0F", X"E5", --5090
  X"CD", X"90", X"11", X"2B", X"CD", X"E5", X"19", X"22", --5098
  X"5B", X"5C", X"FD", X"36", X"07", X"00", X"E1", X"C9", --50A0
  X"FD", X"CB", X"02", X"5E", X"C4", X"1D", X"11", X"A7", --50A8
  X"FD", X"CB", X"01", X"6E", X"C8", X"3A", X"08", X"5C", --50B0
  X"FD", X"CB", X"01", X"AE", X"F5", X"FD", X"CB", X"02", --50B8
  X"6E", X"C4", X"6E", X"0D", X"F1", X"FE", X"20", X"30", --50C0
  X"52", X"FE", X"10", X"30", X"2D", X"FE", X"06", X"30", --50C8
  X"0A", X"47", X"E6", X"01", X"4F", X"78", X"1F", X"C6", --50D0
  X"12", X"18", X"2A", X"20", X"09", X"21", X"6A", X"5C", --50D8
  X"3E", X"08", X"AE", X"77", X"18", X"0E", X"FE", X"0E", --50E0
  X"D8", X"D6", X"0D", X"21", X"41", X"5C", X"BE", X"77", --50E8
  X"20", X"02", X"36", X"00", X"FD", X"CB", X"02", X"DE", --50F0
  X"BF", X"C9", X"47", X"E6", X"07", X"4F", X"3E", X"10", --50F8
  X"CB", X"58", X"20", X"01", X"3C", X"FD", X"71", X"D3", --5100
  X"11", X"0D", X"11", X"18", X"06", X"3A", X"0D", X"5C", --5108
  X"11", X"A8", X"10", X"2A", X"4F", X"5C", X"23", X"23", --5110
  X"73", X"23", X"72", X"37", X"C9", X"CD", X"4D", X"0D", --5118
  X"FD", X"CB", X"02", X"9E", X"FD", X"CB", X"02", X"AE", --5120
  X"2A", X"8A", X"5C", X"E5", X"2A", X"3D", X"5C", X"E5", --5128
  X"21", X"67", X"11", X"E5", X"ED", X"73", X"3D", X"5C", --5130
  X"2A", X"82", X"5C", X"E5", X"37", X"CD", X"95", X"11", --5138
  X"EB", X"CD", X"7D", X"18", X"EB", X"CD", X"E1", X"18", --5140
  X"2A", X"8A", X"5C", X"E3", X"EB", X"CD", X"4D", X"0D", --5148
  X"3A", X"8B", X"5C", X"92", X"38", X"26", X"20", X"06", --5150
  X"7B", X"FD", X"96", X"50", X"30", X"1E", X"3E", X"20", --5158
  X"D5", X"CD", X"F4", X"09", X"D1", X"18", X"E9", X"16", --5160
  X"00", X"FD", X"5E", X"FE", X"21", X"90", X"1A", X"CD", --5168
  X"B5", X"03", X"FD", X"36", X"00", X"FF", X"ED", X"5B", --5170
  X"8A", X"5C", X"18", X"02", X"D1", X"E1", X"E1", X"22", --5178
  X"3D", X"5C", X"C1", X"D5", X"CD", X"D9", X"0D", X"E1", --5180
  X"22", X"82", X"5C", X"FD", X"36", X"26", X"00", X"C9", --5188
  X"2A", X"61", X"5C", X"2B", X"A7", X"ED", X"5B", X"59", --5190
  X"5C", X"FD", X"CB", X"37", X"6E", X"C8", X"ED", X"5B", --5198
  X"61", X"5C", X"D8", X"2A", X"63", X"5C", X"C9", X"7E", --51A0
  X"FE", X"0E", X"01", X"06", X"00", X"CC", X"E8", X"19", --51A8
  X"7E", X"23", X"FE", X"0D", X"20", X"F1", X"C9", X"F3", --51B0
  X"3E", X"FF", X"ED", X"5B", X"B2", X"5C", X"D9", X"ED", --51B8
  X"4B", X"B4", X"5C", X"ED", X"5B", X"38", X"5C", X"2A", --51C0
  X"7B", X"5C", X"D9", X"47", X"3E", X"07", X"D3", X"FE", --51C8
  X"3E", X"3F", X"ED", X"47", X"00", X"00", X"00", X"00", --51D0
  X"00", X"00", X"62", X"6B", X"36", X"02", X"2B", X"BC", --51D8
  X"20", X"FA", X"A7", X"ED", X"52", X"19", X"23", X"30", --51E0
  X"06", X"35", X"28", X"03", X"35", X"28", X"F3", X"2B", --51E8
  X"D9", X"ED", X"43", X"B4", X"5C", X"ED", X"53", X"38", --51F0
  X"5C", X"22", X"7B", X"5C", X"D9", X"04", X"28", X"19", --51F8
  X"22", X"B4", X"5C", X"11", X"AF", X"3E", X"01", X"A8", --5200
  X"00", X"EB", X"ED", X"B8", X"EB", X"23", X"22", X"7B", --5208
  X"5C", X"2B", X"01", X"40", X"00", X"ED", X"43", X"38", --5210
  X"5C", X"22", X"B2", X"5C", X"21", X"00", X"3C", X"22", --5218
  X"36", X"5C", X"2A", X"B2", X"5C", X"36", X"3E", X"2B", --5220
  X"F9", X"2B", X"2B", X"22", X"3D", X"5C", X"ED", X"56", --5228
  X"FD", X"21", X"3A", X"5C", X"FB", X"21", X"B6", X"5C", --5230
  X"22", X"4F", X"5C", X"11", X"AF", X"15", X"01", X"15", --5238
  X"00", X"EB", X"ED", X"B0", X"EB", X"2B", X"22", X"57", --5240
  X"5C", X"23", X"22", X"53", X"5C", X"22", X"4B", X"5C", --5248
  X"36", X"80", X"23", X"22", X"59", X"5C", X"36", X"0D", --5250
  X"23", X"36", X"80", X"23", X"22", X"61", X"5C", X"22", --5258
  X"63", X"5C", X"22", X"65", X"5C", X"3E", X"38", X"32", --5260
  X"8D", X"5C", X"32", X"8F", X"5C", X"32", X"48", X"5C", --5268
  X"21", X"23", X"05", X"22", X"09", X"5C", X"FD", X"35", --5270
  X"C6", X"FD", X"35", X"CA", X"21", X"C6", X"15", X"11", --5278
  X"10", X"5C", X"01", X"0E", X"00", X"ED", X"B0", X"FD", --5280
  X"CB", X"01", X"CE", X"CD", X"DF", X"0E", X"FD", X"36", --5288
  X"31", X"02", X"CD", X"6B", X"0D", X"AF", X"11", X"38", --5290
  X"15", X"CD", X"0A", X"0C", X"FD", X"CB", X"02", X"EE", --5298
  X"18", X"07", X"FD", X"36", X"31", X"02", X"CD", X"95", --52A0
  X"17", X"CD", X"B0", X"16", X"3E", X"00", X"CD", X"01", --52A8
  X"16", X"CD", X"2C", X"0F", X"CD", X"17", X"1B", X"FD", --52B0
  X"CB", X"00", X"7E", X"20", X"12", X"FD", X"CB", X"30", --52B8
  X"66", X"28", X"40", X"2A", X"59", X"5C", X"CD", X"A7", --52C0
  X"11", X"FD", X"36", X"00", X"FF", X"18", X"DD", X"2A", --52C8
  X"59", X"5C", X"22", X"5D", X"5C", X"CD", X"FB", X"19", --52D0
  X"78", X"B1", X"C2", X"5D", X"15", X"DF", X"FE", X"0D", --52D8
  X"28", X"C0", X"FD", X"CB", X"30", X"46", X"C4", X"AF", --52E0
  X"0D", X"CD", X"6E", X"0D", X"3E", X"19", X"FD", X"96", --52E8
  X"4F", X"32", X"8C", X"5C", X"FD", X"CB", X"01", X"FE", --52F0
  X"FD", X"36", X"00", X"FF", X"FD", X"36", X"0A", X"01", --52F8
  X"CD", X"8A", X"1B", X"76", X"FD", X"CB", X"01", X"AE", --5300
  X"FD", X"CB", X"30", X"4E", X"C4", X"CD", X"0E", X"3A", --5308
  X"3A", X"5C", X"3C", X"F5", X"21", X"00", X"00", X"FD", --5310
  X"74", X"37", X"FD", X"74", X"26", X"22", X"0B", X"5C", --5318
  X"21", X"01", X"00", X"22", X"16", X"5C", X"CD", X"B0", --5320
  X"16", X"FD", X"CB", X"37", X"AE", X"CD", X"6E", X"0D", --5328
  X"FD", X"CB", X"02", X"EE", X"F1", X"47", X"FE", X"0A", --5330
  X"38", X"02", X"C6", X"07", X"CD", X"EF", X"15", X"3E", --5338
  X"20", X"D7", X"78", X"11", X"91", X"13", X"CD", X"0A", --5340
  X"0C", X"CD", X"3B", X"3B", X"00", X"CD", X"0A", X"0C", --5348
  X"ED", X"4B", X"45", X"5C", X"CD", X"1B", X"1A", X"3E", --5350
  X"3A", X"D7", X"FD", X"4E", X"0D", X"06", X"00", X"CD", --5358
  X"1B", X"1A", X"CD", X"97", X"10", X"3A", X"3A", X"5C", --5360
  X"3C", X"28", X"1B", X"FE", X"09", X"28", X"04", X"FE", --5368
  X"15", X"20", X"03", X"FD", X"34", X"0D", X"01", X"03", --5370
  X"00", X"11", X"70", X"5C", X"21", X"44", X"5C", X"CB", --5378
  X"7E", X"28", X"01", X"09", X"ED", X"B8", X"FD", X"36", --5380
  X"0A", X"FF", X"FD", X"CB", X"01", X"9E", X"C3", X"AC", --5388
  X"12", X"80", X"4F", X"CB", X"4E", X"45", X"58", X"54", --5390
  X"20", X"77", X"69", X"74", X"68", X"6F", X"75", X"74", --5398
  X"20", X"46", X"4F", X"D2", X"56", X"61", X"72", X"69", --53A0
  X"61", X"62", X"6C", X"65", X"20", X"6E", X"6F", X"74", --53A8
  X"20", X"66", X"6F", X"75", X"6E", X"E4", X"53", X"75", --53B0
  X"62", X"73", X"63", X"72", X"69", X"70", X"74", X"20", --53B8
  X"77", X"72", X"6F", X"6E", X"E7", X"4F", X"75", X"74", --53C0
  X"20", X"6F", X"66", X"20", X"6D", X"65", X"6D", X"6F", --53C8
  X"72", X"F9", X"4F", X"75", X"74", X"20", X"6F", X"66", --53D0
  X"20", X"73", X"63", X"72", X"65", X"65", X"EE", X"4E", --53D8
  X"75", X"6D", X"62", X"65", X"72", X"20", X"74", X"6F", --53E0
  X"6F", X"20", X"62", X"69", X"E7", X"52", X"45", X"54", --53E8
  X"55", X"52", X"4E", X"20", X"77", X"69", X"74", X"68", --53F0
  X"6F", X"75", X"74", X"20", X"47", X"4F", X"53", X"55", --53F8
  X"C2", X"45", X"6E", X"64", X"20", X"6F", X"66", X"20", --5400
  X"66", X"69", X"6C", X"E5", X"53", X"54", X"4F", X"50", --5408
  X"20", X"73", X"74", X"61", X"74", X"65", X"6D", X"65", --5410
  X"6E", X"F4", X"49", X"6E", X"76", X"61", X"6C", X"69", --5418
  X"64", X"20", X"61", X"72", X"67", X"75", X"6D", X"65", --5420
  X"6E", X"F4", X"49", X"6E", X"74", X"65", X"67", X"65", --5428
  X"72", X"20", X"6F", X"75", X"74", X"20", X"6F", X"66", --5430
  X"20", X"72", X"61", X"6E", X"67", X"E5", X"4E", X"6F", --5438
  X"6E", X"73", X"65", X"6E", X"73", X"65", X"20", X"69", --5440
  X"6E", X"20", X"42", X"41", X"53", X"49", X"C3", X"42", --5448
  X"52", X"45", X"41", X"4B", X"20", X"2D", X"20", X"43", --5450
  X"4F", X"4E", X"54", X"20", X"72", X"65", X"70", X"65", --5458
  X"61", X"74", X"F3", X"4F", X"75", X"74", X"20", X"6F", --5460
  X"66", X"20", X"44", X"41", X"54", X"C1", X"49", X"6E", --5468
  X"76", X"61", X"6C", X"69", X"64", X"20", X"66", X"69", --5470
  X"6C", X"65", X"20", X"6E", X"61", X"6D", X"E5", X"4E", --5478
  X"6F", X"20", X"72", X"6F", X"6F", X"6D", X"20", X"66", --5480
  X"6F", X"72", X"20", X"6C", X"69", X"6E", X"E5", X"53", --5488
  X"54", X"4F", X"50", X"20", X"69", X"6E", X"20", X"49", --5490
  X"4E", X"50", X"55", X"D4", X"46", X"4F", X"52", X"20", --5498
  X"77", X"69", X"74", X"68", X"6F", X"75", X"74", X"20", --54A0
  X"4E", X"45", X"58", X"D4", X"49", X"6E", X"76", X"61", --54A8
  X"6C", X"69", X"64", X"20", X"49", X"2F", X"4F", X"20", --54B0
  X"64", X"65", X"76", X"69", X"63", X"E5", X"49", X"6E", --54B8
  X"76", X"61", X"6C", X"69", X"64", X"20", X"63", X"6F", --54C0
  X"6C", X"6F", X"75", X"F2", X"42", X"52", X"45", X"41", --54C8
  X"4B", X"20", X"69", X"6E", X"74", X"6F", X"20", X"70", --54D0
  X"72", X"6F", X"67", X"72", X"61", X"ED", X"52", X"41", --54D8
  X"4D", X"54", X"4F", X"50", X"20", X"6E", X"6F", X"20", --54E0
  X"67", X"6F", X"6F", X"E4", X"53", X"74", X"61", X"74", --54E8
  X"65", X"6D", X"65", X"6E", X"74", X"20", X"6C", X"6F", --54F0
  X"73", X"F4", X"49", X"6E", X"76", X"61", X"6C", X"69", --54F8
  X"64", X"20", X"73", X"74", X"72", X"65", X"61", X"ED", --5500
  X"46", X"4E", X"20", X"77", X"69", X"74", X"68", X"6F", --5508
  X"75", X"74", X"20", X"44", X"45", X"C6", X"50", X"61", --5510
  X"72", X"61", X"6D", X"65", X"74", X"65", X"72", X"20", --5518
  X"65", X"72", X"72", X"6F", X"F2", X"54", X"61", X"70", --5520
  X"65", X"20", X"6C", X"6F", X"61", X"64", X"69", X"6E", --5528
  X"67", X"20", X"65", X"72", X"72", X"6F", X"F2", X"2C", --5530
  X"A0", X"7F", X"20", X"31", X"39", X"38", X"32", X"20", --5538
  X"53", X"69", X"6E", X"63", X"6C", X"61", X"69", X"72", --5540
  X"20", X"52", X"65", X"73", X"65", X"61", X"72", X"63", --5548
  X"68", X"20", X"4C", X"74", X"E4", X"3E", X"10", X"01", --5550
  X"00", X"00", X"C3", X"13", X"13", X"ED", X"43", X"49", --5558
  X"5C", X"2A", X"5D", X"5C", X"EB", X"21", X"55", X"15", --5560
  X"E5", X"2A", X"61", X"5C", X"37", X"ED", X"52", X"E5", --5568
  X"60", X"69", X"CD", X"6E", X"19", X"20", X"06", X"CD", --5570
  X"B8", X"19", X"CD", X"E8", X"19", X"C1", X"79", X"3D", --5578
  X"B0", X"28", X"28", X"C5", X"03", X"03", X"03", X"03", --5580
  X"2B", X"ED", X"5B", X"53", X"5C", X"D5", X"CD", X"55", --5588
  X"16", X"E1", X"22", X"53", X"5C", X"C1", X"C5", X"13", --5590
  X"2A", X"61", X"5C", X"2B", X"2B", X"ED", X"B8", X"2A", --5598
  X"49", X"5C", X"EB", X"C1", X"70", X"2B", X"71", X"2B", --55A0
  X"73", X"2B", X"72", X"F1", X"C3", X"A2", X"12", X"F4", --55A8
  X"09", X"A8", X"10", X"4B", X"F4", X"09", X"C4", X"15", --55B0
  X"53", X"81", X"0F", X"C4", X"15", X"52", X"F4", X"09", --55B8
  X"C4", X"15", X"50", X"80", X"CF", X"12", X"01", X"00", --55C0
  X"06", X"00", X"0B", X"00", X"01", X"00", X"01", X"00", --55C8
  X"06", X"00", X"10", X"00", X"FD", X"CB", X"02", X"6E", --55D0
  X"20", X"04", X"FD", X"CB", X"02", X"DE", X"CD", X"E6", --55D8
  X"15", X"D8", X"28", X"FA", X"CF", X"07", X"D9", X"E5", --55E0
  X"2A", X"51", X"5C", X"23", X"23", X"18", X"08", X"1E", --55E8
  X"30", X"83", X"D9", X"E5", X"2A", X"51", X"5C", X"5E", --55F0
  X"23", X"56", X"EB", X"CD", X"2C", X"16", X"E1", X"D9", --55F8
  X"C9", X"87", X"C6", X"16", X"6F", X"26", X"5C", X"5E", --5600
  X"23", X"56", X"7A", X"B3", X"20", X"02", X"CF", X"17", --5608
  X"1B", X"2A", X"4F", X"5C", X"19", X"22", X"51", X"5C", --5610
  X"FD", X"CB", X"30", X"A6", X"23", X"23", X"23", X"23", --5618
  X"4E", X"21", X"2D", X"16", X"CD", X"DC", X"16", X"D0", --5620
  X"16", X"00", X"5E", X"19", X"E9", X"4B", X"06", X"53", --5628
  X"12", X"50", X"1B", X"00", X"FD", X"CB", X"02", X"C6", --5630
  X"FD", X"CB", X"01", X"AE", X"FD", X"CB", X"30", X"E6", --5638
  X"18", X"04", X"FD", X"CB", X"02", X"86", X"FD", X"CB", --5640
  X"01", X"8E", X"C3", X"4D", X"0D", X"FD", X"CB", X"01", --5648
  X"CE", X"C9", X"01", X"01", X"00", X"E5", X"CD", X"05", --5650
  X"1F", X"E1", X"CD", X"64", X"16", X"2A", X"65", X"5C", --5658
  X"EB", X"ED", X"B8", X"C9", X"F5", X"E5", X"21", X"4B", --5660
  X"5C", X"3E", X"0E", X"5E", X"23", X"56", X"E3", X"A7", --5668
  X"ED", X"52", X"19", X"E3", X"30", X"09", X"D5", X"EB", --5670
  X"09", X"EB", X"72", X"2B", X"73", X"23", X"D1", X"23", --5678
  X"3D", X"20", X"E8", X"EB", X"D1", X"F1", X"A7", X"ED", --5680
  X"52", X"44", X"4D", X"03", X"19", X"EB", X"C9", X"00", --5688
  X"00", X"EB", X"11", X"8F", X"16", X"7E", X"E6", X"C0", --5690
  X"20", X"F7", X"56", X"23", X"5E", X"C9", X"2A", X"63", --5698
  X"5C", X"2B", X"CD", X"55", X"16", X"23", X"23", X"C1", --56A0
  X"ED", X"43", X"61", X"5C", X"C1", X"EB", X"23", X"C9", --56A8
  X"2A", X"59", X"5C", X"36", X"0D", X"22", X"5B", X"5C", --56B0
  X"23", X"36", X"80", X"23", X"22", X"61", X"5C", X"2A", --56B8
  X"61", X"5C", X"22", X"63", X"5C", X"2A", X"63", X"5C", --56C0
  X"22", X"65", X"5C", X"E5", X"21", X"92", X"5C", X"22", --56C8
  X"68", X"5C", X"E1", X"C9", X"ED", X"5B", X"59", X"5C", --56D0
  X"C3", X"E5", X"19", X"23", X"7E", X"A7", X"C8", X"B9", --56D8
  X"23", X"20", X"F8", X"37", X"C9", X"CD", X"1E", X"17", --56E0
  X"CD", X"01", X"17", X"01", X"00", X"00", X"11", X"E2", --56E8
  X"A3", X"EB", X"19", X"38", X"07", X"01", X"D4", X"15", --56F0
  X"09", X"4E", X"23", X"46", X"EB", X"71", X"23", X"70", --56F8
  X"C9", X"E5", X"2A", X"4F", X"5C", X"09", X"23", X"23", --5700
  X"23", X"4E", X"EB", X"21", X"16", X"17", X"CD", X"DC", --5708
  X"16", X"4E", X"06", X"00", X"09", X"E9", X"4B", X"05", --5710
  X"53", X"03", X"50", X"01", X"E1", X"C9", X"CD", X"94", --5718
  X"1E", X"FE", X"10", X"38", X"02", X"CF", X"17", X"C6", --5720
  X"03", X"07", X"21", X"10", X"5C", X"4F", X"06", X"00", --5728
  X"09", X"4E", X"23", X"46", X"2B", X"C9", X"EF", X"01", --5730
  X"38", X"CD", X"1E", X"17", X"78", X"B1", X"28", X"16", --5738
  X"EB", X"2A", X"4F", X"5C", X"09", X"23", X"23", X"23", --5740
  X"7E", X"EB", X"FE", X"4B", X"28", X"08", X"FE", X"53", --5748
  X"28", X"04", X"FE", X"50", X"20", X"CF", X"CD", X"5D", --5750
  X"17", X"73", X"23", X"72", X"C9", X"E5", X"CD", X"F1", --5758
  X"2B", X"78", X"B1", X"20", X"02", X"CF", X"0E", X"C5", --5760
  X"1A", X"E6", X"DF", X"4F", X"21", X"7A", X"17", X"CD", --5768
  X"DC", X"16", X"30", X"F1", X"4E", X"06", X"00", X"09", --5770
  X"C1", X"E9", X"4B", X"06", X"53", X"08", X"50", X"0A", --5778
  X"00", X"1E", X"01", X"18", X"06", X"1E", X"06", X"18", --5780
  X"02", X"1E", X"10", X"0B", X"78", X"B1", X"20", X"D5", --5788
  X"57", X"E1", X"C9", X"18", X"90", X"ED", X"73", X"3F", --5790
  X"5C", X"FD", X"36", X"02", X"10", X"CD", X"AF", X"0D", --5798
  X"FD", X"CB", X"02", X"C6", X"FD", X"46", X"31", X"CD", --57A0
  X"44", X"0E", X"FD", X"CB", X"02", X"86", X"FD", X"CB", --57A8
  X"30", X"C6", X"2A", X"49", X"5C", X"ED", X"5B", X"6C", --57B0
  X"5C", X"A7", X"ED", X"52", X"19", X"38", X"22", X"D5", --57B8
  X"CD", X"6E", X"19", X"11", X"C0", X"02", X"EB", X"ED", --57C0
  X"52", X"E3", X"CD", X"6E", X"19", X"C1", X"C5", X"CD", --57C8
  X"B8", X"19", X"C1", X"09", X"38", X"0E", X"EB", X"56", --57D0
  X"23", X"5E", X"2B", X"ED", X"53", X"6C", X"5C", X"18", --57D8
  X"ED", X"22", X"6C", X"5C", X"2A", X"6C", X"5C", X"CD", --57E0
  X"6E", X"19", X"28", X"01", X"EB", X"CD", X"33", X"18", --57E8
  X"FD", X"CB", X"02", X"A6", X"C9", X"3E", X"03", X"18", --57F0
  X"02", X"3E", X"02", X"FD", X"36", X"02", X"00", X"CD", --57F8
  X"30", X"25", X"C4", X"01", X"16", X"DF", X"CD", X"70", --5800
  X"20", X"38", X"14", X"DF", X"FE", X"3B", X"28", X"04", --5808
  X"FE", X"2C", X"20", X"06", X"E7", X"CD", X"82", X"1C", --5810
  X"18", X"08", X"CD", X"E6", X"1C", X"18", X"03", X"CD", --5818
  X"DE", X"1C", X"CD", X"EE", X"1B", X"CD", X"99", X"1E", --5820
  X"78", X"E6", X"3F", X"67", X"69", X"22", X"49", X"5C", --5828
  X"CD", X"6E", X"19", X"1E", X"01", X"CD", X"55", X"18", --5830
  X"D7", X"FD", X"CB", X"02", X"66", X"28", X"F6", X"3A", --5838
  X"6B", X"5C", X"FD", X"96", X"4F", X"20", X"EE", X"AB", --5840
  X"C8", X"E5", X"D5", X"21", X"6C", X"5C", X"CD", X"0F", --5848
  X"19", X"D1", X"E1", X"18", X"E0", X"ED", X"4B", X"49", --5850
  X"5C", X"CD", X"80", X"19", X"16", X"3E", X"28", X"05", --5858
  X"11", X"00", X"00", X"CB", X"13", X"FD", X"73", X"2D", --5860
  X"7E", X"FE", X"40", X"C1", X"D0", X"C5", X"CD", X"28", --5868
  X"1A", X"23", X"23", X"23", X"FD", X"CB", X"01", X"86", --5870
  X"7A", X"A7", X"28", X"05", X"D7", X"FD", X"CB", X"01", --5878
  X"C6", X"D5", X"EB", X"FD", X"CB", X"30", X"96", X"21", --5880
  X"3B", X"5C", X"CB", X"96", X"FD", X"CB", X"37", X"6E", --5888
  X"28", X"02", X"CB", X"D6", X"2A", X"5F", X"5C", X"A7", --5890
  X"ED", X"52", X"20", X"05", X"3E", X"3F", X"CD", X"C1", --5898
  X"18", X"CD", X"E1", X"18", X"EB", X"7E", X"CD", X"B6", --58A0
  X"18", X"23", X"FE", X"0D", X"28", X"06", X"EB", X"CD", --58A8
  X"37", X"19", X"18", X"E0", X"D1", X"C9", X"FE", X"0E", --58B0
  X"C0", X"23", X"23", X"23", X"23", X"23", X"23", X"7E", --58B8
  X"C9", X"D9", X"2A", X"8F", X"5C", X"E5", X"CB", X"BC", --58C0
  X"CB", X"FD", X"22", X"8F", X"5C", X"21", X"91", X"5C", --58C8
  X"56", X"D5", X"36", X"00", X"CD", X"F4", X"09", X"E1", --58D0
  X"FD", X"74", X"57", X"E1", X"22", X"8F", X"5C", X"D9", --58D8
  X"C9", X"2A", X"5B", X"5C", X"A7", X"ED", X"52", X"C0", --58E0
  X"3A", X"41", X"5C", X"CB", X"07", X"28", X"04", X"C6", --58E8
  X"43", X"18", X"16", X"21", X"3B", X"5C", X"CB", X"9E", --58F0
  X"3E", X"4B", X"CB", X"56", X"28", X"0B", X"CB", X"DE", --58F8
  X"3C", X"FD", X"CB", X"30", X"5E", X"28", X"02", X"3E", --5900
  X"43", X"D5", X"CD", X"C1", X"18", X"D1", X"C9", X"5E", --5908
  X"23", X"56", X"E5", X"EB", X"23", X"CD", X"6E", X"19", --5910
  X"CD", X"95", X"16", X"E1", X"FD", X"CB", X"37", X"6E", --5918
  X"C0", X"72", X"2B", X"73", X"C9", X"7B", X"A7", X"F8", --5920
  X"18", X"0D", X"AF", X"09", X"3C", X"38", X"FC", X"ED", --5928
  X"42", X"3D", X"28", X"F1", X"C3", X"EF", X"15", X"CD", --5930
  X"1B", X"2D", X"30", X"30", X"FE", X"21", X"38", X"2C", --5938
  X"FD", X"CB", X"01", X"96", X"FE", X"CB", X"28", X"24", --5940
  X"FE", X"3A", X"20", X"0E", X"FD", X"CB", X"37", X"6E", --5948
  X"20", X"16", X"FD", X"CB", X"30", X"56", X"28", X"14", --5950
  X"18", X"0E", X"FE", X"22", X"20", X"0A", X"F5", X"3A", --5958
  X"6A", X"5C", X"EE", X"04", X"32", X"6A", X"5C", X"F1", --5960
  X"FD", X"CB", X"01", X"D6", X"D7", X"C9", X"E5", X"2A", --5968
  X"53", X"5C", X"54", X"5D", X"C1", X"CD", X"80", X"19", --5970
  X"D0", X"C5", X"CD", X"B8", X"19", X"EB", X"18", X"F4", --5978
  X"7E", X"B8", X"C0", X"23", X"7E", X"2B", X"B9", X"C9", --5980
  X"23", X"23", X"23", X"22", X"5D", X"5C", X"0E", X"00", --5988
  X"15", X"C8", X"E7", X"BB", X"20", X"04", X"A7", X"C9", --5990
  X"23", X"7E", X"CD", X"B6", X"18", X"22", X"5D", X"5C", --5998
  X"FE", X"22", X"20", X"01", X"0D", X"FE", X"3A", X"28", --59A0
  X"04", X"FE", X"CB", X"20", X"04", X"CB", X"41", X"28", --59A8
  X"DF", X"FE", X"0D", X"20", X"E3", X"15", X"37", X"C9", --59B0
  X"E5", X"7E", X"FE", X"40", X"38", X"17", X"CB", X"6F", --59B8
  X"28", X"14", X"87", X"FA", X"C7", X"19", X"3F", X"01", --59C0
  X"05", X"00", X"30", X"02", X"0E", X"12", X"17", X"23", --59C8
  X"7E", X"30", X"FB", X"18", X"06", X"23", X"23", X"4E", --59D0
  X"23", X"46", X"23", X"09", X"D1", X"A7", X"ED", X"52", --59D8
  X"44", X"4D", X"19", X"EB", X"C9", X"CD", X"DD", X"19", --59E0
  X"C5", X"78", X"2F", X"47", X"79", X"2F", X"4F", X"03", --59E8
  X"CD", X"64", X"16", X"EB", X"E1", X"19", X"D5", X"ED", --59F0
  X"B0", X"E1", X"C9", X"2A", X"59", X"5C", X"2B", X"22", --59F8
  X"5D", X"5C", X"E7", X"21", X"92", X"5C", X"22", X"65", --5A00
  X"5C", X"CD", X"3B", X"2D", X"CD", X"A2", X"2D", X"38", --5A08
  X"04", X"21", X"F0", X"D8", X"09", X"DA", X"8A", X"1C", --5A10
  X"C3", X"C5", X"16", X"D5", X"E5", X"AF", X"CB", X"78", --5A18
  X"20", X"20", X"60", X"69", X"1E", X"FF", X"18", X"08", --5A20
  X"D5", X"56", X"23", X"5E", X"E5", X"EB", X"1E", X"20", --5A28
  X"01", X"18", X"FC", X"CD", X"2A", X"19", X"01", X"9C", --5A30
  X"FF", X"CD", X"2A", X"19", X"0E", X"F6", X"CD", X"2A", --5A38
  X"19", X"7D", X"CD", X"EF", X"15", X"E1", X"D1", X"C9", --5A40
  X"B1", X"CB", X"BC", X"BF", X"C4", X"AF", X"B4", X"93", --5A48
  X"91", X"92", X"95", X"98", X"98", X"98", X"98", X"98", --5A50
  X"98", X"98", X"7F", X"81", X"2E", X"6C", X"6E", X"70", --5A58
  X"48", X"94", X"56", X"3F", X"41", X"2B", X"17", X"1F", --5A60
  X"37", X"77", X"44", X"0F", X"59", X"2B", X"43", X"2D", --5A68
  X"51", X"3A", X"6D", X"42", X"0D", X"49", X"5C", X"44", --5A70
  X"15", X"5D", X"01", X"3D", X"02", X"06", X"00", X"67", --5A78
  X"1E", X"06", X"CB", X"05", X"F0", X"1C", X"06", X"00", --5A80
  X"ED", X"1E", X"00", X"EE", X"1C", X"00", X"23", X"1F", --5A88
  X"04", X"3D", X"06", X"CC", X"06", X"05", X"03", X"1D", --5A90
  X"04", X"00", X"AB", X"1D", X"05", X"CD", X"1F", X"05", --5A98
  X"89", X"20", X"05", X"02", X"2C", X"05", X"B2", X"1B", --5AA0
  X"00", X"B7", X"11", X"03", X"A1", X"1E", X"05", X"F9", --5AA8
  X"17", X"08", X"00", X"80", X"1E", X"03", X"4F", X"1E", --5AB0
  X"00", X"5F", X"1E", X"03", X"AC", X"1E", X"00", X"6B", --5AB8
  X"0D", X"09", X"00", X"DC", X"22", X"06", X"00", X"3A", --5AC0
  X"1F", X"05", X"ED", X"1D", X"05", X"27", X"1E", X"03", --5AC8
  X"42", X"1E", X"09", X"05", X"82", X"23", X"00", X"AC", --5AD0
  X"0E", X"05", X"C9", X"1F", X"05", X"F5", X"17", X"0B", --5AD8
  X"0B", X"0B", X"0B", X"08", X"00", X"F8", X"03", X"09", --5AE0
  X"05", X"20", X"23", X"07", X"07", X"07", X"07", X"07", --5AE8
  X"07", X"08", X"00", X"7A", X"1E", X"06", X"00", X"94", --5AF0
  X"22", X"05", X"60", X"1F", X"06", X"2C", X"0A", X"00", --5AF8
  X"36", X"17", X"06", X"00", X"E5", X"16", X"0A", X"00", --5B00
  X"93", X"17", X"0A", X"2C", X"0A", X"00", X"93", X"17", --5B08
  X"0A", X"00", X"93", X"17", X"00", X"93", X"17", X"FD", --5B10
  X"CB", X"01", X"BE", X"CD", X"FB", X"19", X"AF", X"32", --5B18
  X"47", X"5C", X"3D", X"32", X"3A", X"5C", X"18", X"01", --5B20
  X"E7", X"CD", X"BF", X"16", X"FD", X"34", X"0D", X"FA", --5B28
  X"8A", X"1C", X"DF", X"06", X"00", X"FE", X"0D", X"28", --5B30
  X"7A", X"FE", X"3A", X"28", X"EB", X"21", X"76", X"1B", --5B38
  X"E5", X"4F", X"E7", X"79", X"D6", X"CE", X"DA", X"8A", --5B40
  X"1C", X"4F", X"21", X"48", X"1A", X"09", X"4E", X"09", --5B48
  X"18", X"03", X"2A", X"74", X"5C", X"7E", X"23", X"22", --5B50
  X"74", X"5C", X"01", X"52", X"1B", X"C5", X"4F", X"FE", --5B58
  X"20", X"30", X"0C", X"21", X"01", X"1C", X"06", X"00", --5B60
  X"09", X"4E", X"09", X"E5", X"DF", X"05", X"C9", X"DF", --5B68
  X"B9", X"C2", X"8A", X"1C", X"E7", X"C9", X"CD", X"54", --5B70
  X"1F", X"38", X"02", X"CF", X"14", X"CD", X"4D", X"3B", --5B78
  X"00", X"20", X"71", X"2A", X"42", X"5C", X"CB", X"7C", --5B80
  X"28", X"14", X"21", X"FE", X"FF", X"22", X"45", X"5C", --5B88
  X"2A", X"61", X"5C", X"2B", X"ED", X"5B", X"59", X"5C", --5B90
  X"1B", X"3A", X"44", X"5C", X"18", X"33", X"CD", X"6E", --5B98
  X"19", X"3A", X"44", X"5C", X"28", X"19", X"A7", X"20", --5BA0
  X"43", X"47", X"7E", X"E6", X"C0", X"78", X"28", X"0F", --5BA8
  X"CF", X"FF", X"C1", X"CD", X"30", X"25", X"C8", X"2A", --5BB0
  X"55", X"5C", X"3E", X"C0", X"A6", X"C0", X"AF", X"FE", --5BB8
  X"01", X"CE", X"00", X"56", X"23", X"5E", X"ED", X"53", --5BC0
  X"45", X"5C", X"23", X"5E", X"23", X"56", X"EB", X"19", --5BC8
  X"23", X"22", X"55", X"5C", X"EB", X"22", X"5D", X"5C", --5BD0
  X"57", X"1E", X"00", X"FD", X"36", X"0A", X"FF", X"15", --5BD8
  X"FD", X"72", X"0D", X"CA", X"28", X"1B", X"14", X"CD", --5BE0
  X"8B", X"19", X"28", X"08", X"CF", X"16", X"CD", X"30", --5BE8
  X"25", X"C0", X"C1", X"C1", X"CD", X"5D", X"3B", X"28", --5BF0
  X"BA", X"FE", X"3A", X"CA", X"28", X"1B", X"C3", X"8A", --5BF8
  X"1C", X"0F", X"1D", X"4B", X"09", X"67", X"0B", X"7B", --5C00
  X"8E", X"71", X"B4", X"81", X"CF", X"CD", X"DE", X"1C", --5C08
  X"BF", X"C1", X"CC", X"EE", X"1B", X"EB", X"2A", X"74", --5C10
  X"5C", X"4E", X"23", X"46", X"EB", X"C5", X"C9", X"CD", --5C18
  X"B2", X"28", X"FD", X"36", X"37", X"00", X"30", X"08", --5C20
  X"FD", X"CB", X"37", X"CE", X"20", X"18", X"CF", X"01", --5C28
  X"CC", X"96", X"29", X"FD", X"CB", X"01", X"76", X"20", --5C30
  X"0D", X"AF", X"CD", X"30", X"25", X"C4", X"F1", X"2B", --5C38
  X"21", X"71", X"5C", X"B6", X"77", X"EB", X"ED", X"43", --5C40
  X"72", X"5C", X"22", X"4D", X"5C", X"C9", X"C1", X"CD", --5C48
  X"56", X"1C", X"CD", X"EE", X"1B", X"C9", X"3A", X"3B", --5C50
  X"5C", X"F5", X"CD", X"FB", X"24", X"F1", X"FD", X"56", --5C58
  X"01", X"AA", X"E6", X"40", X"20", X"24", X"CB", X"7A", --5C60
  X"C2", X"FF", X"2A", X"C9", X"CD", X"B2", X"28", X"F5", --5C68
  X"79", X"F6", X"9F", X"3C", X"20", X"14", X"F1", X"18", --5C70
  X"A9", X"E7", X"CD", X"82", X"1C", X"FE", X"2C", X"20", --5C78
  X"09", X"E7", X"CD", X"FB", X"24", X"FD", X"CB", X"01", --5C80
  X"76", X"C0", X"CF", X"0B", X"CD", X"FB", X"24", X"FD", --5C88
  X"CB", X"01", X"76", X"C8", X"18", X"F4", X"FD", X"CB", --5C90
  X"01", X"7E", X"FD", X"CB", X"02", X"86", X"C4", X"4D", --5C98
  X"0D", X"F1", X"3A", X"74", X"5C", X"D6", X"13", X"CD", --5CA0
  X"FC", X"21", X"CD", X"EE", X"1B", X"2A", X"8F", X"5C", --5CA8
  X"22", X"8D", X"5C", X"21", X"91", X"5C", X"7E", X"07", --5CB0
  X"AE", X"E6", X"AA", X"AE", X"77", X"C9", X"CD", X"30", --5CB8
  X"25", X"28", X"13", X"FD", X"CB", X"02", X"86", X"CD", --5CC0
  X"4D", X"0D", X"21", X"90", X"5C", X"7E", X"F6", X"F8", --5CC8
  X"77", X"FD", X"CB", X"57", X"B6", X"DF", X"CD", X"E2", --5CD0
  X"21", X"18", X"9F", X"C3", X"05", X"06", X"FE", X"0D", --5CD8
  X"28", X"04", X"FE", X"3A", X"20", X"9C", X"CD", X"30", --5CE0
  X"25", X"C8", X"EF", X"A0", X"38", X"C9", X"CF", X"08", --5CE8
  X"C1", X"CD", X"30", X"25", X"28", X"0A", X"EF", X"02", --5CF0
  X"38", X"EB", X"CD", X"E9", X"34", X"DA", X"B3", X"1B", --5CF8
  X"C3", X"29", X"1B", X"FE", X"CD", X"20", X"09", X"E7", --5D00
  X"CD", X"82", X"1C", X"CD", X"EE", X"1B", X"18", X"06", --5D08
  X"CD", X"EE", X"1B", X"EF", X"A1", X"38", X"EF", X"C0", --5D10
  X"02", X"01", X"E0", X"01", X"38", X"CD", X"FF", X"2A", --5D18
  X"22", X"68", X"5C", X"2B", X"7E", X"CB", X"FE", X"01", --5D20
  X"06", X"00", X"09", X"07", X"38", X"06", X"0E", X"0D", --5D28
  X"CD", X"55", X"16", X"23", X"E5", X"EF", X"02", X"02", --5D30
  X"38", X"E1", X"EB", X"0E", X"0A", X"ED", X"B0", X"2A", --5D38
  X"45", X"5C", X"EB", X"73", X"23", X"72", X"FD", X"56", --5D40
  X"0D", X"14", X"23", X"72", X"CD", X"DA", X"1D", X"D0", --5D48
  X"FD", X"46", X"38", X"2A", X"45", X"5C", X"22", X"42", --5D50
  X"5C", X"3A", X"47", X"5C", X"ED", X"44", X"57", X"2A", --5D58
  X"5D", X"5C", X"1E", X"F3", X"C5", X"ED", X"4B", X"55", --5D60
  X"5C", X"CD", X"86", X"1D", X"ED", X"43", X"55", X"5C", --5D68
  X"C1", X"38", X"11", X"E7", X"F6", X"20", X"B8", X"28", --5D70
  X"03", X"E7", X"18", X"E8", X"E7", X"3E", X"01", X"92", --5D78
  X"32", X"44", X"5C", X"C9", X"CF", X"11", X"7E", X"FE", --5D80
  X"3A", X"28", X"18", X"23", X"7E", X"E6", X"C0", X"37", --5D88
  X"C0", X"46", X"23", X"4E", X"ED", X"43", X"42", X"5C", --5D90
  X"23", X"4E", X"23", X"46", X"E5", X"09", X"44", X"4D", --5D98
  X"E1", X"16", X"00", X"C5", X"CD", X"8B", X"19", X"C1", --5DA0
  X"D0", X"18", X"E0", X"FD", X"CB", X"37", X"4E", X"C2", --5DA8
  X"2E", X"1C", X"2A", X"4D", X"5C", X"CB", X"7E", X"28", --5DB0
  X"1F", X"23", X"22", X"68", X"5C", X"EF", X"E0", X"E2", --5DB8
  X"0F", X"C0", X"02", X"38", X"CD", X"DA", X"1D", X"D8", --5DC0
  X"2A", X"68", X"5C", X"11", X"0F", X"00", X"19", X"5E", --5DC8
  X"23", X"56", X"23", X"66", X"EB", X"C3", X"73", X"1E", --5DD0
  X"CF", X"00", X"EF", X"E1", X"E0", X"E2", X"36", X"00", --5DD8
  X"02", X"01", X"03", X"37", X"00", X"04", X"38", X"A7", --5DE0
  X"C9", X"38", X"37", X"C9", X"E7", X"CD", X"1F", X"1C", --5DE8
  X"CD", X"30", X"25", X"28", X"29", X"DF", X"22", X"5F", --5DF0
  X"5C", X"2A", X"57", X"5C", X"7E", X"FE", X"2C", X"28", --5DF8
  X"09", X"1E", X"E4", X"CD", X"86", X"1D", X"30", X"02", --5E00
  X"CF", X"0D", X"CD", X"77", X"00", X"CD", X"56", X"1C", --5E08
  X"DF", X"22", X"57", X"5C", X"2A", X"5F", X"5C", X"FD", --5E10
  X"36", X"26", X"00", X"CD", X"78", X"00", X"DF", X"FE", --5E18
  X"2C", X"28", X"C9", X"CD", X"EE", X"1B", X"C9", X"CD", --5E20
  X"30", X"25", X"20", X"0B", X"CD", X"FB", X"24", X"FE", --5E28
  X"2C", X"C4", X"EE", X"1B", X"E7", X"18", X"F5", X"3E", --5E30
  X"E4", X"47", X"ED", X"B9", X"11", X"00", X"02", X"C3", --5E38
  X"8B", X"19", X"CD", X"99", X"1E", X"60", X"69", X"CD", --5E40
  X"6E", X"19", X"2B", X"22", X"57", X"5C", X"C9", X"CD", --5E48
  X"99", X"1E", X"78", X"B1", X"20", X"04", X"ED", X"4B", --5E50
  X"78", X"5C", X"ED", X"43", X"76", X"5C", X"C9", X"2A", --5E58
  X"6E", X"5C", X"FD", X"56", X"36", X"18", X"0C", X"CD", --5E60
  X"99", X"1E", X"60", X"69", X"16", X"00", X"7C", X"FE", --5E68
  X"F0", X"30", X"2C", X"22", X"42", X"5C", X"FD", X"72", --5E70
  X"0A", X"C9", X"CD", X"85", X"1E", X"ED", X"79", X"C9", --5E78
  X"CD", X"85", X"1E", X"02", X"C9", X"CD", X"D5", X"2D", --5E80
  X"38", X"15", X"28", X"02", X"ED", X"44", X"F5", X"CD", --5E88
  X"99", X"1E", X"F1", X"C9", X"CD", X"D5", X"2D", X"18", --5E90
  X"03", X"CD", X"A2", X"2D", X"38", X"01", X"C8", X"CF", --5E98
  X"0A", X"CD", X"67", X"1E", X"01", X"00", X"00", X"CD", --5EA0
  X"45", X"1E", X"18", X"03", X"CD", X"99", X"1E", X"78", --5EA8
  X"B1", X"20", X"04", X"ED", X"4B", X"B2", X"5C", X"C5", --5EB0
  X"ED", X"5B", X"4B", X"5C", X"2A", X"59", X"5C", X"2B", --5EB8
  X"CD", X"E5", X"19", X"CD", X"6B", X"0D", X"2A", X"65", --5EC0
  X"5C", X"11", X"32", X"00", X"19", X"D1", X"ED", X"52", --5EC8
  X"30", X"08", X"2A", X"B4", X"5C", X"A7", X"ED", X"52", --5ED0
  X"30", X"02", X"CF", X"15", X"EB", X"22", X"B2", X"5C", --5ED8
  X"D1", X"C1", X"36", X"3E", X"2B", X"F9", X"C5", X"ED", --5EE0
  X"73", X"3D", X"5C", X"EB", X"E9", X"D1", X"FD", X"66", --5EE8
  X"0D", X"24", X"E3", X"33", X"ED", X"4B", X"45", X"5C", --5EF0
  X"C5", X"E5", X"ED", X"73", X"3D", X"5C", X"D5", X"CD", --5EF8
  X"67", X"1E", X"01", X"14", X"00", X"2A", X"65", X"5C", --5F00
  X"09", X"38", X"0A", X"EB", X"21", X"50", X"00", X"19", --5F08
  X"38", X"03", X"ED", X"72", X"D8", X"2E", X"03", X"C3", --5F10
  X"55", X"00", X"01", X"00", X"00", X"CD", X"05", X"1F", --5F18
  X"44", X"4D", X"C9", X"C1", X"E1", X"D1", X"7A", X"FE", --5F20
  X"3E", X"28", X"0B", X"3B", X"E3", X"EB", X"ED", X"73", --5F28
  X"3D", X"5C", X"C5", X"C3", X"73", X"1E", X"D5", X"E5", --5F30
  X"CF", X"06", X"CD", X"99", X"1E", X"76", X"0B", X"78", --5F38
  X"B1", X"28", X"0C", X"78", X"A1", X"3C", X"20", X"01", --5F40
  X"03", X"FD", X"CB", X"01", X"6E", X"28", X"EE", X"FD", --5F48
  X"CB", X"01", X"AE", X"C9", X"3E", X"7F", X"DB", X"FE", --5F50
  X"1F", X"D8", X"3E", X"FE", X"DB", X"FE", X"1F", X"C9", --5F58
  X"CD", X"30", X"25", X"28", X"05", X"3E", X"CE", X"C3", --5F60
  X"39", X"1E", X"FD", X"CB", X"01", X"F6", X"CD", X"8D", --5F68
  X"2C", X"30", X"16", X"E7", X"FE", X"24", X"20", X"05", --5F70
  X"FD", X"CB", X"01", X"B6", X"E7", X"FE", X"28", X"20", --5F78
  X"3C", X"E7", X"FE", X"29", X"28", X"20", X"CD", X"8D", --5F80
  X"2C", X"D2", X"8A", X"1C", X"EB", X"E7", X"FE", X"24", --5F88
  X"20", X"02", X"EB", X"E7", X"EB", X"01", X"06", X"00", --5F90
  X"CD", X"55", X"16", X"23", X"23", X"36", X"0E", X"FE", --5F98
  X"2C", X"20", X"03", X"E7", X"18", X"E0", X"FE", X"29", --5FA0
  X"20", X"13", X"E7", X"FE", X"3D", X"20", X"0E", X"E7", --5FA8
  X"3A", X"3B", X"5C", X"F5", X"CD", X"FB", X"24", X"F1", --5FB0
  X"FD", X"AE", X"01", X"E6", X"40", X"C2", X"8A", X"1C", --5FB8
  X"CD", X"EE", X"1B", X"CD", X"30", X"25", X"E1", X"C8", --5FC0
  X"E9", X"3E", X"03", X"18", X"02", X"3E", X"02", X"CD", --5FC8
  X"30", X"25", X"C4", X"01", X"16", X"CD", X"4D", X"0D", --5FD0
  X"CD", X"DF", X"1F", X"CD", X"EE", X"1B", X"C9", X"DF", --5FD8
  X"CD", X"45", X"20", X"28", X"0D", X"CD", X"4E", X"20", --5FE0
  X"28", X"FB", X"CD", X"FC", X"1F", X"CD", X"4E", X"20", --5FE8
  X"28", X"F3", X"FE", X"29", X"C8", X"CD", X"C3", X"1F", --5FF0
  X"3E", X"0D", X"D7", X"C9", X"DF", X"FE", X"AC", X"20", --5FF8
  X"0D", X"CD", X"79", X"1C", X"CD", X"C3", X"1F", X"CD", --6000
  X"07", X"23", X"3E", X"16", X"18", X"10", X"FE", X"AD", --6008
  X"20", X"12", X"E7", X"CD", X"82", X"1C", X"CD", X"C3", --6010
  X"1F", X"CD", X"99", X"1E", X"3E", X"17", X"D7", X"79", --6018
  X"D7", X"78", X"D7", X"C9", X"CD", X"F2", X"21", X"D0", --6020
  X"CD", X"70", X"20", X"D0", X"CD", X"FB", X"24", X"CD", --6028
  X"C3", X"1F", X"FD", X"CB", X"01", X"76", X"CC", X"F1", --6030
  X"2B", X"C2", X"E3", X"2D", X"78", X"B1", X"0B", X"C8", --6038
  X"1A", X"13", X"D7", X"18", X"F7", X"FE", X"29", X"C8", --6040
  X"FE", X"0D", X"C8", X"FE", X"3A", X"C9", X"DF", X"FE", --6048
  X"3B", X"28", X"14", X"FE", X"2C", X"20", X"0A", X"CD", --6050
  X"30", X"25", X"28", X"0B", X"3E", X"06", X"D7", X"18", --6058
  X"06", X"FE", X"27", X"C0", X"CD", X"F5", X"1F", X"E7", --6060
  X"CD", X"45", X"20", X"20", X"01", X"C1", X"BF", X"C9", --6068
  X"FE", X"23", X"37", X"C0", X"E7", X"CD", X"82", X"1C", --6070
  X"A7", X"CD", X"C3", X"1F", X"CD", X"94", X"1E", X"FE", --6078
  X"10", X"D2", X"0E", X"16", X"CD", X"01", X"16", X"A7", --6080
  X"C9", X"CD", X"30", X"25", X"28", X"08", X"3E", X"01", --6088
  X"CD", X"01", X"16", X"CD", X"6E", X"0D", X"FD", X"36", --6090
  X"02", X"01", X"CD", X"C1", X"20", X"CD", X"EE", X"1B", --6098
  X"ED", X"4B", X"88", X"5C", X"3A", X"6B", X"5C", X"B8", --60A0
  X"38", X"03", X"0E", X"21", X"47", X"ED", X"43", X"88", --60A8
  X"5C", X"3E", X"19", X"90", X"32", X"8C", X"5C", X"FD", --60B0
  X"CB", X"02", X"86", X"CD", X"D9", X"0D", X"C3", X"6E", --60B8
  X"0D", X"CD", X"4E", X"20", X"28", X"FB", X"FE", X"28", --60C0
  X"20", X"0E", X"E7", X"CD", X"DF", X"1F", X"DF", X"FE", --60C8
  X"29", X"C2", X"8A", X"1C", X"E7", X"C3", X"B2", X"21", --60D0
  X"FE", X"CA", X"20", X"11", X"E7", X"CD", X"1F", X"1C", --60D8
  X"FD", X"CB", X"37", X"FE", X"FD", X"CB", X"01", X"76", --60E0
  X"C2", X"8A", X"1C", X"18", X"0D", X"CD", X"8D", X"2C", --60E8
  X"D2", X"AF", X"21", X"CD", X"1F", X"1C", X"FD", X"CB", --60F0
  X"37", X"BE", X"CD", X"30", X"25", X"CA", X"B2", X"21", --60F8
  X"CD", X"BF", X"16", X"21", X"71", X"5C", X"CB", X"B6", --6100
  X"CB", X"EE", X"01", X"01", X"00", X"CB", X"7E", X"20", --6108
  X"0B", X"3A", X"3B", X"5C", X"E6", X"40", X"20", X"02", --6110
  X"0E", X"03", X"B6", X"77", X"F7", X"36", X"0D", X"79", --6118
  X"0F", X"0F", X"30", X"05", X"3E", X"22", X"12", X"2B", --6120
  X"77", X"22", X"5B", X"5C", X"FD", X"CB", X"37", X"7E", --6128
  X"20", X"2C", X"2A", X"5D", X"5C", X"E5", X"2A", X"3D", --6130
  X"5C", X"E5", X"21", X"3A", X"21", X"E5", X"FD", X"CB", --6138
  X"30", X"66", X"28", X"04", X"ED", X"73", X"3D", X"5C", --6140
  X"2A", X"61", X"5C", X"CD", X"A7", X"11", X"FD", X"36", --6148
  X"00", X"FF", X"CD", X"2C", X"0F", X"FD", X"CB", X"01", --6150
  X"BE", X"CD", X"B9", X"21", X"18", X"03", X"CD", X"2C", --6158
  X"0F", X"FD", X"36", X"22", X"00", X"CD", X"D6", X"21", --6160
  X"20", X"0A", X"CD", X"1D", X"11", X"ED", X"4B", X"82", --6168
  X"5C", X"CD", X"D9", X"0D", X"21", X"71", X"5C", X"CB", --6170
  X"AE", X"CB", X"7E", X"CB", X"BE", X"20", X"1C", X"E1", --6178
  X"E1", X"22", X"3D", X"5C", X"E1", X"22", X"5F", X"5C", --6180
  X"FD", X"CB", X"01", X"FE", X"CD", X"B9", X"21", X"2A", --6188
  X"5F", X"5C", X"FD", X"36", X"26", X"00", X"22", X"5D", --6190
  X"5C", X"18", X"17", X"2A", X"63", X"5C", X"ED", X"5B", --6198
  X"61", X"5C", X"37", X"ED", X"52", X"44", X"4D", X"CD", --61A0
  X"B2", X"2A", X"CD", X"FF", X"2A", X"18", X"03", X"CD", --61A8
  X"FC", X"1F", X"CD", X"4E", X"20", X"CA", X"C1", X"20", --61B0
  X"C9", X"2A", X"61", X"5C", X"22", X"5D", X"5C", X"DF", --61B8
  X"FE", X"E2", X"28", X"0C", X"3A", X"71", X"5C", X"CD", --61C0
  X"59", X"1C", X"DF", X"FE", X"0D", X"C8", X"CF", X"0B", --61C8
  X"CD", X"30", X"25", X"C8", X"CF", X"10", X"2A", X"51", --61D0
  X"5C", X"23", X"23", X"23", X"23", X"7E", X"FE", X"4B", --61D8
  X"C9", X"E7", X"CD", X"F2", X"21", X"D8", X"DF", X"FE", --61E0
  X"2C", X"28", X"F6", X"FE", X"3B", X"28", X"F2", X"C3", --61E8
  X"8A", X"1C", X"FE", X"D9", X"D8", X"FE", X"DF", X"3F", --61F0
  X"D8", X"F5", X"E7", X"F1", X"D6", X"C9", X"F5", X"CD", --61F8
  X"82", X"1C", X"F1", X"A7", X"CD", X"C3", X"1F", X"F5", --6200
  X"CD", X"94", X"1E", X"57", X"F1", X"D7", X"7A", X"D7", --6208
  X"C9", X"D6", X"11", X"CE", X"00", X"28", X"1D", X"D6", --6210
  X"02", X"CE", X"00", X"28", X"56", X"FE", X"01", X"7A", --6218
  X"06", X"01", X"20", X"04", X"07", X"07", X"06", X"04", --6220
  X"4F", X"7A", X"FE", X"02", X"30", X"16", X"79", X"21", --6228
  X"91", X"5C", X"18", X"38", X"7A", X"06", X"07", X"38", --6230
  X"05", X"07", X"07", X"07", X"06", X"38", X"4F", X"7A", --6238
  X"FE", X"0A", X"38", X"02", X"CF", X"13", X"21", X"8F", --6240
  X"5C", X"FE", X"08", X"38", X"0B", X"7E", X"28", X"07", --6248
  X"B0", X"2F", X"E6", X"24", X"28", X"01", X"78", X"4F", --6250
  X"79", X"CD", X"6C", X"22", X"3E", X"07", X"BA", X"9F", --6258
  X"CD", X"6C", X"22", X"07", X"07", X"E6", X"50", X"47", --6260
  X"3E", X"08", X"BA", X"9F", X"AE", X"A0", X"AE", X"77", --6268
  X"23", X"78", X"C9", X"9F", X"7A", X"0F", X"06", X"80", --6270
  X"20", X"03", X"0F", X"06", X"40", X"4F", X"7A", X"FE", --6278
  X"08", X"28", X"04", X"FE", X"02", X"30", X"BD", X"79", --6280
  X"21", X"8F", X"5C", X"CD", X"6C", X"22", X"79", X"0F", --6288
  X"0F", X"0F", X"18", X"D8", X"CD", X"94", X"1E", X"FE", --6290
  X"08", X"30", X"A9", X"D3", X"FE", X"07", X"07", X"07", --6298
  X"CB", X"6F", X"20", X"02", X"EE", X"07", X"32", X"48", --62A0
  X"5C", X"C9", X"3E", X"AF", X"90", X"DA", X"F9", X"24", --62A8
  X"47", X"A7", X"1F", X"37", X"1F", X"A7", X"1F", X"A8", --62B0
  X"E6", X"F8", X"A8", X"67", X"79", X"07", X"07", X"07", --62B8
  X"A8", X"E6", X"C7", X"A8", X"07", X"07", X"6F", X"79", --62C0
  X"E6", X"07", X"C9", X"CD", X"07", X"23", X"CD", X"AA", --62C8
  X"22", X"47", X"04", X"7E", X"07", X"10", X"FD", X"E6", --62D0
  X"01", X"C3", X"28", X"2D", X"CD", X"07", X"23", X"CD", --62D8
  X"E5", X"22", X"C3", X"4D", X"0D", X"ED", X"43", X"7D", --62E0
  X"5C", X"CD", X"AA", X"22", X"47", X"04", X"3E", X"FE", --62E8
  X"0F", X"10", X"FD", X"47", X"7E", X"FD", X"4E", X"57", --62F0
  X"CB", X"41", X"20", X"01", X"A0", X"CB", X"51", X"20", --62F8
  X"02", X"A8", X"2F", X"77", X"C3", X"DB", X"0B", X"CD", --6300
  X"14", X"23", X"47", X"C5", X"CD", X"14", X"23", X"59", --6308
  X"C1", X"51", X"4F", X"C9", X"CD", X"D5", X"2D", X"DA", --6310
  X"F9", X"24", X"0E", X"01", X"C8", X"0E", X"FF", X"C9", --6318
  X"DF", X"FE", X"2C", X"C2", X"8A", X"1C", X"E7", X"CD", --6320
  X"82", X"1C", X"CD", X"EE", X"1B", X"EF", X"2A", X"3D", --6328
  X"38", X"7E", X"FE", X"81", X"30", X"05", X"EF", X"02", --6330
  X"38", X"18", X"A1", X"EF", X"A3", X"38", X"36", X"83", --6338
  X"EF", X"C5", X"02", X"38", X"CD", X"7D", X"24", X"C5", --6340
  X"EF", X"31", X"E1", X"04", X"38", X"7E", X"FE", X"80", --6348
  X"30", X"08", X"EF", X"02", X"02", X"38", X"C1", X"C3", --6350
  X"DC", X"22", X"EF", X"C2", X"01", X"C0", X"02", X"03", --6358
  X"01", X"E0", X"0F", X"C0", X"01", X"31", X"E0", X"01", --6360
  X"31", X"E0", X"A0", X"C1", X"02", X"38", X"FD", X"34", --6368
  X"62", X"CD", X"94", X"1E", X"6F", X"E5", X"CD", X"94", --6370
  X"1E", X"E1", X"67", X"22", X"7D", X"5C", X"C1", X"C3", --6378
  X"20", X"24", X"DF", X"FE", X"2C", X"28", X"06", X"CD", --6380
  X"EE", X"1B", X"C3", X"77", X"24", X"E7", X"CD", X"82", --6388
  X"1C", X"CD", X"EE", X"1B", X"EF", X"C5", X"A2", X"04", --6390
  X"1F", X"31", X"30", X"30", X"00", X"06", X"02", X"38", --6398
  X"C3", X"77", X"24", X"C0", X"02", X"C1", X"02", X"31", --63A0
  X"2A", X"E1", X"01", X"E1", X"2A", X"0F", X"E0", X"05", --63A8
  X"2A", X"E0", X"01", X"3D", X"38", X"7E", X"FE", X"81", --63B0
  X"30", X"07", X"EF", X"02", X"02", X"38", X"C3", X"77", --63B8
  X"24", X"CD", X"7D", X"24", X"C5", X"EF", X"02", X"E1", --63C0
  X"01", X"05", X"C1", X"02", X"01", X"31", X"E1", X"04", --63C8
  X"C2", X"02", X"01", X"31", X"E1", X"04", X"E2", X"E5", --63D0
  X"E0", X"03", X"A2", X"04", X"31", X"1F", X"C5", X"02", --63D8
  X"20", X"C0", X"02", X"C2", X"02", X"C1", X"E5", X"04", --63E0
  X"E0", X"E2", X"04", X"0F", X"E1", X"01", X"C1", X"02", --63E8
  X"E0", X"04", X"E2", X"E5", X"04", X"03", X"C2", X"2A", --63F0
  X"E1", X"2A", X"0F", X"02", X"38", X"1A", X"FE", X"81", --63F8
  X"C1", X"DA", X"77", X"24", X"C5", X"EF", X"01", X"38", --6400
  X"3A", X"7D", X"5C", X"CD", X"28", X"2D", X"EF", X"C0", --6408
  X"0F", X"01", X"38", X"3A", X"7E", X"5C", X"CD", X"28", --6410
  X"2D", X"EF", X"C5", X"0F", X"E0", X"E5", X"38", X"C1", --6418
  X"05", X"28", X"3C", X"18", X"14", X"EF", X"E1", X"31", --6420
  X"E3", X"04", X"E2", X"E4", X"04", X"03", X"C1", X"02", --6428
  X"E4", X"04", X"E2", X"E3", X"04", X"0F", X"C2", X"02", --6430
  X"38", X"C5", X"EF", X"C0", X"02", X"E1", X"0F", X"31", --6438
  X"38", X"3A", X"7D", X"5C", X"CD", X"28", X"2D", X"EF", --6440
  X"03", X"E0", X"E2", X"0F", X"C0", X"01", X"E0", X"38", --6448
  X"3A", X"7E", X"5C", X"CD", X"28", X"2D", X"EF", X"03", --6450
  X"38", X"CD", X"B7", X"24", X"C1", X"10", X"C6", X"EF", --6458
  X"02", X"02", X"01", X"38", X"3A", X"7D", X"5C", X"CD", --6460
  X"28", X"2D", X"EF", X"03", X"01", X"38", X"3A", X"7E", --6468
  X"5C", X"CD", X"28", X"2D", X"EF", X"03", X"38", X"CD", --6470
  X"B7", X"24", X"C3", X"4D", X"0D", X"EF", X"31", X"28", --6478
  X"34", X"32", X"00", X"01", X"05", X"E5", X"01", X"05", --6480
  X"2A", X"38", X"CD", X"D5", X"2D", X"38", X"06", X"E6", --6488
  X"FC", X"C6", X"04", X"30", X"02", X"3E", X"FC", X"F5", --6490
  X"CD", X"28", X"2D", X"EF", X"E5", X"01", X"05", X"31", --6498
  X"1F", X"C4", X"02", X"31", X"A2", X"04", X"1F", X"C1", --64A0
  X"01", X"C0", X"02", X"31", X"04", X"31", X"0F", X"A1", --64A8
  X"03", X"1B", X"C3", X"02", X"38", X"C1", X"C9", X"CD", --64B0
  X"07", X"23", X"79", X"B8", X"30", X"06", X"69", X"D5", --64B8
  X"AF", X"5F", X"18", X"07", X"B1", X"C8", X"68", X"41", --64C0
  X"D5", X"16", X"00", X"60", X"78", X"1F", X"85", X"38", --64C8
  X"03", X"BC", X"38", X"07", X"94", X"4F", X"D9", X"C1", --64D0
  X"C5", X"18", X"04", X"4F", X"D5", X"D9", X"C1", X"2A", --64D8
  X"7D", X"5C", X"78", X"84", X"47", X"79", X"3C", X"85", --64E0
  X"38", X"0D", X"28", X"0D", X"3D", X"4F", X"CD", X"E5", --64E8
  X"22", X"D9", X"79", X"10", X"D9", X"D1", X"C9", X"28", --64F0
  X"F3", X"CF", X"0A", X"DF", X"06", X"00", X"C5", X"4F", --64F8
  X"21", X"96", X"25", X"CD", X"DC", X"16", X"79", X"D2", --6500
  X"84", X"26", X"06", X"00", X"4E", X"09", X"E9", X"CD", --6508
  X"74", X"00", X"03", X"FE", X"0D", X"CA", X"8A", X"1C", --6510
  X"FE", X"22", X"20", X"F3", X"CD", X"74", X"00", X"FE", --6518
  X"22", X"C9", X"E7", X"FE", X"28", X"20", X"06", X"CD", --6520
  X"79", X"1C", X"DF", X"FE", X"29", X"C2", X"8A", X"1C", --6528
  X"FD", X"CB", X"01", X"7E", X"C9", X"CD", X"07", X"23", --6530
  X"2A", X"36", X"5C", X"11", X"00", X"01", X"19", X"79", --6538
  X"0F", X"0F", X"0F", X"E6", X"E0", X"A8", X"5F", X"79", --6540
  X"E6", X"18", X"EE", X"40", X"57", X"06", X"60", X"C5", --6548
  X"D5", X"E5", X"1A", X"AE", X"28", X"04", X"3C", X"20", --6550
  X"1A", X"3D", X"4F", X"06", X"07", X"14", X"23", X"1A", --6558
  X"AE", X"A9", X"20", X"0F", X"10", X"F7", X"C1", X"C1", --6560
  X"C1", X"3E", X"80", X"90", X"01", X"01", X"00", X"F7", --6568
  X"12", X"18", X"0A", X"E1", X"11", X"08", X"00", X"19", --6570
  X"D1", X"C1", X"10", X"D3", X"48", X"C3", X"B2", X"2A", --6578
  X"CD", X"07", X"23", X"79", X"0F", X"0F", X"0F", X"4F", --6580
  X"E6", X"E0", X"A8", X"6F", X"79", X"E6", X"03", X"EE", --6588
  X"58", X"67", X"7E", X"C3", X"28", X"2D", X"22", X"1C", --6590
  X"28", X"4F", X"2E", X"F2", X"2B", X"12", X"A8", X"56", --6598
  X"A5", X"57", X"A7", X"84", X"A6", X"8F", X"C4", X"E6", --65A0
  X"AA", X"BF", X"AB", X"C7", X"A9", X"CE", X"00", X"E7", --65A8
  X"C3", X"FF", X"24", X"DF", X"23", X"E5", X"01", X"00", --65B0
  X"00", X"CD", X"0F", X"25", X"20", X"1B", X"CD", X"0F", --65B8
  X"25", X"28", X"FB", X"CD", X"30", X"25", X"28", X"11", --65C0
  X"F7", X"E1", X"D5", X"7E", X"23", X"12", X"13", X"FE", --65C8
  X"22", X"20", X"F8", X"7E", X"23", X"FE", X"22", X"28", --65D0
  X"F2", X"0B", X"D1", X"21", X"3B", X"5C", X"CB", X"B6", --65D8
  X"CB", X"7E", X"C4", X"B2", X"2A", X"C3", X"12", X"27", --65E0
  X"E7", X"CD", X"FB", X"24", X"FE", X"29", X"C2", X"8A", --65E8
  X"1C", X"E7", X"C3", X"12", X"27", X"C3", X"BD", X"27", --65F0
  X"CD", X"30", X"25", X"28", X"28", X"ED", X"4B", X"76", --65F8
  X"5C", X"CD", X"2B", X"2D", X"EF", X"A1", X"0F", X"34", --6600
  X"37", X"16", X"04", X"34", X"80", X"41", X"00", X"00", --6608
  X"80", X"32", X"02", X"A1", X"03", X"31", X"38", X"CD", --6610
  X"A2", X"2D", X"ED", X"43", X"76", X"5C", X"7E", X"A7", --6618
  X"28", X"03", X"D6", X"10", X"77", X"18", X"09", X"CD", --6620
  X"30", X"25", X"28", X"04", X"EF", X"A3", X"38", X"34", --6628
  X"E7", X"C3", X"C3", X"26", X"01", X"5A", X"10", X"E7", --6630
  X"FE", X"23", X"CA", X"0D", X"27", X"21", X"3B", X"5C", --6638
  X"CB", X"B6", X"CB", X"7E", X"28", X"1F", X"C3", X"6C", --6640
  X"3B", X"0E", X"00", X"20", X"13", X"CD", X"1E", X"03", --6648
  X"30", X"0E", X"15", X"5F", X"CD", X"33", X"03", X"F5", --6650
  X"01", X"01", X"00", X"F7", X"F1", X"12", X"0E", X"01", --6658
  X"06", X"00", X"CD", X"B2", X"2A", X"C3", X"12", X"27", --6660
  X"CD", X"22", X"25", X"C4", X"35", X"25", X"E7", X"C3", --6668
  X"DB", X"25", X"CD", X"22", X"25", X"C4", X"80", X"25", --6670
  X"E7", X"18", X"48", X"CD", X"22", X"25", X"C4", X"CB", --6678
  X"22", X"E7", X"18", X"3F", X"CD", X"88", X"2C", X"30", --6680
  X"56", X"FE", X"41", X"30", X"3C", X"CD", X"30", X"25", --6688
  X"20", X"23", X"CD", X"9B", X"2C", X"DF", X"01", X"06", --6690
  X"00", X"CD", X"55", X"16", X"23", X"36", X"0E", X"23", --6698
  X"EB", X"2A", X"65", X"5C", X"0E", X"05", X"A7", X"ED", --66A0
  X"42", X"22", X"65", X"5C", X"ED", X"B0", X"EB", X"2B", --66A8
  X"CD", X"77", X"00", X"18", X"0E", X"DF", X"23", X"7E", --66B0
  X"FE", X"0E", X"20", X"FA", X"23", X"CD", X"B4", X"33", --66B8
  X"22", X"5D", X"5C", X"FD", X"CB", X"01", X"F6", X"18", --66C0
  X"14", X"CD", X"B2", X"28", X"DA", X"2E", X"1C", X"CC", --66C8
  X"96", X"29", X"3A", X"3B", X"5C", X"FE", X"C0", X"38", --66D0
  X"04", X"23", X"CD", X"B4", X"33", X"18", X"33", X"01", --66D8
  X"DB", X"09", X"FE", X"2D", X"28", X"27", X"01", X"18", --66E0
  X"10", X"FE", X"AE", X"28", X"20", X"D6", X"AF", X"DA", --66E8
  X"8A", X"1C", X"01", X"F0", X"04", X"FE", X"14", X"28", --66F0
  X"14", X"D2", X"8A", X"1C", X"06", X"10", X"C6", X"DC", --66F8
  X"4F", X"FE", X"DF", X"30", X"02", X"CB", X"B1", X"FE", --6700
  X"EE", X"38", X"02", X"CB", X"B9", X"C5", X"E7", X"C3", --6708
  X"FF", X"24", X"DF", X"FE", X"28", X"20", X"0C", X"FD", --6710
  X"CB", X"01", X"76", X"20", X"17", X"CD", X"52", X"2A", --6718
  X"E7", X"18", X"F0", X"06", X"00", X"4F", X"21", X"95", --6720
  X"27", X"CD", X"DC", X"16", X"30", X"06", X"4E", X"21", --6728
  X"ED", X"26", X"09", X"46", X"D1", X"7A", X"B8", X"38", --6730
  X"3A", X"A7", X"CA", X"18", X"00", X"C5", X"21", X"3B", --6738
  X"5C", X"7B", X"FE", X"ED", X"20", X"06", X"CB", X"76", --6740
  X"20", X"02", X"1E", X"99", X"D5", X"CD", X"30", X"25", --6748
  X"28", X"09", X"7B", X"E6", X"3F", X"47", X"EF", X"3B", --6750
  X"38", X"18", X"09", X"7B", X"FD", X"AE", X"01", X"E6", --6758
  X"40", X"C2", X"8A", X"1C", X"D1", X"21", X"3B", X"5C", --6760
  X"CB", X"F6", X"CB", X"7B", X"20", X"02", X"CB", X"B6", --6768
  X"C1", X"18", X"C1", X"D5", X"79", X"FD", X"CB", X"01", --6770
  X"76", X"20", X"15", X"E6", X"3F", X"C6", X"08", X"4F", --6778
  X"FE", X"10", X"20", X"04", X"CB", X"F1", X"18", X"08", --6780
  X"38", X"D7", X"FE", X"17", X"28", X"02", X"CB", X"F9", --6788
  X"C5", X"E7", X"C3", X"FF", X"24", X"2B", X"CF", X"2D", --6790
  X"C3", X"2A", X"C4", X"2F", X"C5", X"5E", X"C6", X"3D", --6798
  X"CE", X"3E", X"CC", X"3C", X"CD", X"C7", X"C9", X"C8", --67A0
  X"CA", X"C9", X"CB", X"C5", X"C7", X"C6", X"C8", X"00", --67A8
  X"06", X"08", X"08", X"0A", X"02", X"03", X"05", X"05", --67B0
  X"05", X"05", X"05", X"05", X"06", X"CD", X"30", X"25", --67B8
  X"20", X"35", X"E7", X"CD", X"8D", X"2C", X"D2", X"8A", --67C0
  X"1C", X"E7", X"FE", X"24", X"F5", X"20", X"01", X"E7", --67C8
  X"FE", X"28", X"20", X"12", X"E7", X"FE", X"29", X"28", --67D0
  X"10", X"CD", X"FB", X"24", X"DF", X"FE", X"2C", X"20", --67D8
  X"03", X"E7", X"18", X"F5", X"FE", X"29", X"C2", X"8A", --67E0
  X"1C", X"E7", X"21", X"3B", X"5C", X"CB", X"B6", X"F1", --67E8
  X"28", X"02", X"CB", X"F6", X"C3", X"12", X"27", X"E7", --67F0
  X"E6", X"DF", X"47", X"E7", X"D6", X"24", X"4F", X"20", --67F8
  X"01", X"E7", X"E7", X"E5", X"2A", X"53", X"5C", X"2B", --6800
  X"11", X"CE", X"00", X"C5", X"CD", X"86", X"1D", X"C1", --6808
  X"30", X"02", X"CF", X"18", X"E5", X"CD", X"AB", X"28", --6810
  X"E6", X"DF", X"B8", X"20", X"08", X"CD", X"AB", X"28", --6818
  X"D6", X"24", X"B9", X"28", X"0C", X"E1", X"2B", X"11", --6820
  X"00", X"02", X"C5", X"CD", X"8B", X"19", X"C1", X"18", --6828
  X"D7", X"A7", X"CC", X"AB", X"28", X"D1", X"D1", X"ED", --6830
  X"53", X"5D", X"5C", X"CD", X"AB", X"28", X"E5", X"FE", --6838
  X"29", X"28", X"42", X"23", X"7E", X"FE", X"0E", X"16", --6840
  X"40", X"28", X"07", X"2B", X"CD", X"AB", X"28", X"23", --6848
  X"16", X"00", X"23", X"E5", X"D5", X"CD", X"FB", X"24", --6850
  X"F1", X"FD", X"AE", X"01", X"E6", X"40", X"20", X"2B", --6858
  X"E1", X"EB", X"2A", X"65", X"5C", X"01", X"05", X"00", --6860
  X"ED", X"42", X"22", X"65", X"5C", X"ED", X"B0", X"EB", --6868
  X"2B", X"CD", X"AB", X"28", X"FE", X"29", X"28", X"0D", --6870
  X"E5", X"DF", X"FE", X"2C", X"20", X"0D", X"E7", X"E1", --6878
  X"CD", X"AB", X"28", X"18", X"BE", X"E5", X"DF", X"FE", --6880
  X"29", X"28", X"02", X"CF", X"19", X"D1", X"EB", X"22", --6888
  X"5D", X"5C", X"2A", X"0B", X"5C", X"E3", X"22", X"0B", --6890
  X"5C", X"D5", X"E7", X"E7", X"CD", X"FB", X"24", X"E1", --6898
  X"22", X"5D", X"5C", X"E1", X"22", X"0B", X"5C", X"E7", --68A0
  X"C3", X"12", X"27", X"23", X"7E", X"FE", X"21", X"38", --68A8
  X"FA", X"C9", X"FD", X"CB", X"01", X"F6", X"DF", X"CD", --68B0
  X"8D", X"2C", X"D2", X"8A", X"1C", X"E5", X"E6", X"1F", --68B8
  X"4F", X"E7", X"E5", X"FE", X"28", X"28", X"28", X"CB", --68C0
  X"F1", X"FE", X"24", X"28", X"11", X"CB", X"E9", X"CD", --68C8
  X"88", X"2C", X"30", X"0F", X"CD", X"88", X"2C", X"30", --68D0
  X"16", X"CB", X"B1", X"E7", X"18", X"F6", X"E7", X"FD", --68D8
  X"CB", X"01", X"B6", X"3A", X"0C", X"5C", X"A7", X"28", --68E0
  X"06", X"CD", X"30", X"25", X"C2", X"51", X"29", X"41", --68E8
  X"CD", X"30", X"25", X"20", X"08", X"79", X"E6", X"E0", --68F0
  X"CB", X"FF", X"4F", X"18", X"37", X"2A", X"4B", X"5C", --68F8
  X"7E", X"E6", X"7F", X"28", X"2D", X"B9", X"20", X"22", --6900
  X"17", X"87", X"F2", X"3F", X"29", X"38", X"30", X"D1", --6908
  X"D5", X"E5", X"23", X"1A", X"13", X"FE", X"20", X"28", --6910
  X"FA", X"F6", X"20", X"BE", X"28", X"F4", X"F6", X"80", --6918
  X"BE", X"20", X"06", X"1A", X"CD", X"88", X"2C", X"30", --6920
  X"15", X"E1", X"C5", X"CD", X"B8", X"19", X"EB", X"C1", --6928
  X"18", X"CE", X"CB", X"F8", X"D1", X"DF", X"FE", X"28", --6930
  X"28", X"09", X"CB", X"E8", X"18", X"0D", X"D1", X"D1", --6938
  X"D1", X"E5", X"DF", X"CD", X"88", X"2C", X"30", X"03", --6940
  X"E7", X"18", X"F8", X"E1", X"CB", X"10", X"CB", X"70", --6948
  X"C9", X"2A", X"0B", X"5C", X"7E", X"FE", X"29", X"CA", --6950
  X"EF", X"28", X"7E", X"F6", X"60", X"47", X"23", X"7E", --6958
  X"FE", X"0E", X"28", X"07", X"2B", X"CD", X"AB", X"28", --6960
  X"23", X"CB", X"A8", X"78", X"B9", X"28", X"12", X"23", --6968
  X"23", X"23", X"23", X"23", X"CD", X"AB", X"28", X"FE", --6970
  X"29", X"CA", X"EF", X"28", X"CD", X"AB", X"28", X"18", --6978
  X"D9", X"CB", X"69", X"20", X"0C", X"23", X"ED", X"5B", --6980
  X"65", X"5C", X"CD", X"C0", X"33", X"EB", X"22", X"65", --6988
  X"5C", X"D1", X"D1", X"AF", X"3C", X"C9", X"AF", X"47", --6990
  X"CB", X"79", X"20", X"4B", X"CB", X"7E", X"20", X"0E", --6998
  X"3C", X"23", X"4E", X"23", X"46", X"23", X"EB", X"CD", --69A0
  X"B2", X"2A", X"DF", X"C3", X"49", X"2A", X"23", X"23", --69A8
  X"23", X"46", X"CB", X"71", X"28", X"0A", X"05", X"28", --69B0
  X"E8", X"EB", X"DF", X"FE", X"28", X"20", X"61", X"EB", --69B8
  X"EB", X"18", X"24", X"E5", X"DF", X"E1", X"FE", X"2C", --69C0
  X"28", X"20", X"CB", X"79", X"28", X"52", X"CB", X"71", --69C8
  X"20", X"06", X"FE", X"29", X"20", X"3C", X"E7", X"C9", --69D0
  X"FE", X"29", X"28", X"6C", X"FE", X"CC", X"20", X"32", --69D8
  X"DF", X"2B", X"22", X"5D", X"5C", X"18", X"5E", X"21", --69E0
  X"00", X"00", X"E5", X"E7", X"E1", X"79", X"FE", X"C0", --69E8
  X"20", X"09", X"DF", X"FE", X"29", X"28", X"51", X"FE", --69F0
  X"CC", X"28", X"E5", X"C5", X"E5", X"CD", X"EE", X"2A", --69F8
  X"E3", X"EB", X"CD", X"CC", X"2A", X"38", X"19", X"0B", --6A00
  X"CD", X"F4", X"2A", X"09", X"D1", X"C1", X"10", X"B3", --6A08
  X"CB", X"79", X"20", X"66", X"E5", X"CB", X"71", X"20", --6A10
  X"13", X"42", X"4B", X"DF", X"FE", X"29", X"28", X"02", --6A18
  X"CF", X"02", X"E7", X"E1", X"11", X"05", X"00", X"CD", --6A20
  X"F4", X"2A", X"09", X"C9", X"CD", X"EE", X"2A", X"E3", --6A28
  X"CD", X"F4", X"2A", X"C1", X"09", X"23", X"42", X"4B", --6A30
  X"EB", X"CD", X"B1", X"2A", X"DF", X"FE", X"29", X"28", --6A38
  X"07", X"FE", X"2C", X"20", X"DB", X"CD", X"52", X"2A", --6A40
  X"E7", X"FE", X"28", X"28", X"F8", X"FD", X"CB", X"01", --6A48
  X"B6", X"C9", X"CD", X"30", X"25", X"C4", X"F1", X"2B", --6A50
  X"E7", X"FE", X"29", X"28", X"50", X"D5", X"AF", X"F5", --6A58
  X"C5", X"11", X"01", X"00", X"DF", X"E1", X"FE", X"CC", --6A60
  X"28", X"17", X"F1", X"CD", X"CD", X"2A", X"F5", X"50", --6A68
  X"59", X"E5", X"DF", X"E1", X"FE", X"CC", X"28", X"09", --6A70
  X"FE", X"29", X"C2", X"8A", X"1C", X"62", X"6B", X"18", --6A78
  X"13", X"E5", X"E7", X"E1", X"FE", X"29", X"28", X"0C", --6A80
  X"F1", X"CD", X"CD", X"2A", X"F5", X"DF", X"60", X"69", --6A88
  X"FE", X"29", X"20", X"E6", X"F1", X"E3", X"19", X"2B", --6A90
  X"E3", X"A7", X"ED", X"52", X"01", X"00", X"00", X"38", --6A98
  X"07", X"23", X"A7", X"FA", X"20", X"2A", X"44", X"4D", --6AA0
  X"D1", X"FD", X"CB", X"01", X"B6", X"CD", X"30", X"25", --6AA8
  X"C8", X"AF", X"FD", X"CB", X"01", X"B6", X"C5", X"CD", --6AB0
  X"A9", X"33", X"C1", X"2A", X"65", X"5C", X"77", X"23", --6AB8
  X"73", X"23", X"72", X"23", X"71", X"23", X"70", X"23", --6AC0
  X"22", X"65", X"5C", X"C9", X"AF", X"D5", X"E5", X"F5", --6AC8
  X"CD", X"82", X"1C", X"F1", X"CD", X"30", X"25", X"28", --6AD0
  X"12", X"F5", X"CD", X"99", X"1E", X"D1", X"78", X"B1", --6AD8
  X"37", X"28", X"05", X"E1", X"E5", X"A7", X"ED", X"42", --6AE0
  X"7A", X"DE", X"00", X"E1", X"D1", X"C9", X"EB", X"23", --6AE8
  X"5E", X"23", X"56", X"C9", X"CD", X"30", X"25", X"C8", --6AF0
  X"CD", X"A9", X"30", X"DA", X"15", X"1F", X"C9", X"2A", --6AF8
  X"4D", X"5C", X"FD", X"CB", X"37", X"4E", X"28", X"5E", --6B00
  X"01", X"05", X"00", X"03", X"23", X"7E", X"FE", X"20", --6B08
  X"28", X"FA", X"30", X"0B", X"FE", X"10", X"38", X"11", --6B10
  X"FE", X"16", X"30", X"0D", X"23", X"18", X"ED", X"CD", --6B18
  X"88", X"2C", X"38", X"E7", X"FE", X"24", X"CA", X"C0", --6B20
  X"2B", X"79", X"2A", X"59", X"5C", X"2B", X"CD", X"55", --6B28
  X"16", X"23", X"23", X"EB", X"D5", X"2A", X"4D", X"5C", --6B30
  X"1B", X"D6", X"06", X"47", X"28", X"11", X"23", X"7E", --6B38
  X"FE", X"21", X"38", X"FA", X"F6", X"20", X"13", X"12", --6B40
  X"10", X"F4", X"F6", X"80", X"12", X"3E", X"C0", X"2A", --6B48
  X"4D", X"5C", X"AE", X"F6", X"20", X"E1", X"CD", X"EA", --6B50
  X"2B", X"E5", X"EF", X"02", X"38", X"E1", X"01", X"05", --6B58
  X"00", X"A7", X"ED", X"42", X"18", X"40", X"FD", X"CB", --6B60
  X"01", X"76", X"28", X"06", X"11", X"06", X"00", X"19", --6B68
  X"18", X"E7", X"2A", X"4D", X"5C", X"ED", X"4B", X"72", --6B70
  X"5C", X"FD", X"CB", X"37", X"46", X"20", X"30", X"78", --6B78
  X"B1", X"C8", X"E5", X"F7", X"D5", X"C5", X"54", X"5D", --6B80
  X"23", X"36", X"20", X"ED", X"B8", X"E5", X"CD", X"F1", --6B88
  X"2B", X"E1", X"E3", X"A7", X"ED", X"42", X"09", X"30", --6B90
  X"02", X"44", X"4D", X"E3", X"EB", X"78", X"B1", X"28", --6B98
  X"02", X"ED", X"B0", X"C1", X"D1", X"E1", X"EB", X"78", --6BA0
  X"B1", X"C8", X"D5", X"ED", X"B0", X"E1", X"C9", X"2B", --6BA8
  X"2B", X"2B", X"7E", X"E5", X"C5", X"CD", X"C6", X"2B", --6BB0
  X"C1", X"E1", X"03", X"03", X"03", X"C3", X"E8", X"19", --6BB8
  X"3E", X"DF", X"2A", X"4D", X"5C", X"A6", X"F5", X"CD", --6BC0
  X"F1", X"2B", X"EB", X"09", X"C5", X"2B", X"22", X"4D", --6BC8
  X"5C", X"03", X"03", X"03", X"2A", X"59", X"5C", X"2B", --6BD0
  X"CD", X"55", X"16", X"2A", X"4D", X"5C", X"C1", X"C5", --6BD8
  X"03", X"ED", X"B8", X"EB", X"23", X"C1", X"70", X"2B", --6BE0
  X"71", X"F1", X"2B", X"77", X"2A", X"59", X"5C", X"2B", --6BE8
  X"C9", X"2A", X"65", X"5C", X"2B", X"46", X"2B", X"4E", --6BF0
  X"2B", X"56", X"2B", X"5E", X"2B", X"7E", X"22", X"65", --6BF8
  X"5C", X"C9", X"CD", X"B2", X"28", X"C2", X"8A", X"1C", --6C00
  X"CD", X"30", X"25", X"20", X"08", X"CB", X"B1", X"CD", --6C08
  X"96", X"29", X"CD", X"EE", X"1B", X"38", X"08", X"C5", --6C10
  X"CD", X"B8", X"19", X"CD", X"E8", X"19", X"C1", X"CB", --6C18
  X"F9", X"06", X"00", X"C5", X"21", X"01", X"00", X"CB", --6C20
  X"71", X"20", X"02", X"2E", X"05", X"EB", X"E7", X"26", --6C28
  X"FF", X"CD", X"CC", X"2A", X"DA", X"20", X"2A", X"E1", --6C30
  X"C5", X"24", X"E5", X"60", X"69", X"CD", X"F4", X"2A", --6C38
  X"EB", X"DF", X"FE", X"2C", X"28", X"E8", X"FE", X"29", --6C40
  X"20", X"BB", X"E7", X"C1", X"79", X"68", X"26", X"00", --6C48
  X"23", X"23", X"29", X"19", X"DA", X"15", X"1F", X"D5", --6C50
  X"C5", X"E5", X"44", X"4D", X"2A", X"59", X"5C", X"2B", --6C58
  X"CD", X"55", X"16", X"23", X"77", X"C1", X"0B", X"0B", --6C60
  X"0B", X"23", X"71", X"23", X"70", X"C1", X"78", X"23", --6C68
  X"77", X"62", X"6B", X"1B", X"36", X"00", X"CB", X"71", --6C70
  X"28", X"02", X"36", X"20", X"C1", X"ED", X"B8", X"C1", --6C78
  X"70", X"2B", X"71", X"2B", X"3D", X"20", X"F8", X"C9", --6C80
  X"CD", X"1B", X"2D", X"3F", X"D8", X"FE", X"41", X"3F", --6C88
  X"D0", X"FE", X"5B", X"D8", X"FE", X"61", X"3F", X"D0", --6C90
  X"FE", X"7B", X"C9", X"FE", X"C4", X"20", X"19", X"11", --6C98
  X"00", X"00", X"E7", X"D6", X"31", X"CE", X"00", X"20", --6CA0
  X"0A", X"EB", X"3F", X"ED", X"6A", X"DA", X"AD", X"31", --6CA8
  X"EB", X"18", X"EF", X"42", X"4B", X"C3", X"2B", X"2D", --6CB0
  X"FE", X"2E", X"28", X"0F", X"CD", X"3B", X"2D", X"FE", --6CB8
  X"2E", X"20", X"28", X"E7", X"CD", X"1B", X"2D", X"38", --6CC0
  X"22", X"18", X"0A", X"E7", X"CD", X"1B", X"2D", X"DA", --6CC8
  X"8A", X"1C", X"EF", X"A0", X"38", X"EF", X"A1", X"C0", --6CD0
  X"02", X"38", X"DF", X"CD", X"22", X"2D", X"38", X"0B", --6CD8
  X"EF", X"E0", X"A4", X"05", X"C0", X"04", X"0F", X"38", --6CE0
  X"E7", X"18", X"EF", X"FE", X"45", X"28", X"03", X"FE", --6CE8
  X"65", X"C0", X"06", X"FF", X"E7", X"FE", X"2B", X"28", --6CF0
  X"05", X"FE", X"2D", X"20", X"02", X"04", X"E7", X"CD", --6CF8
  X"1B", X"2D", X"38", X"CB", X"C5", X"CD", X"3B", X"2D", --6D00
  X"CD", X"D5", X"2D", X"C1", X"DA", X"AD", X"31", X"A7", --6D08
  X"FA", X"AD", X"31", X"04", X"28", X"02", X"ED", X"44", --6D10
  X"C3", X"4F", X"2D", X"FE", X"30", X"D8", X"FE", X"3A", --6D18
  X"3F", X"C9", X"CD", X"1B", X"2D", X"D8", X"D6", X"30", --6D20
  X"4F", X"06", X"00", X"FD", X"21", X"3A", X"5C", X"AF", --6D28
  X"5F", X"51", X"48", X"47", X"CD", X"B6", X"2A", X"EF", --6D30
  X"38", X"A7", X"C9", X"F5", X"EF", X"A0", X"38", X"F1", --6D38
  X"CD", X"22", X"2D", X"D8", X"EF", X"01", X"A4", X"04", --6D40
  X"0F", X"38", X"CD", X"74", X"00", X"18", X"F1", X"07", --6D48
  X"0F", X"30", X"02", X"2F", X"3C", X"F5", X"21", X"92", --6D50
  X"5C", X"CD", X"0B", X"35", X"EF", X"A4", X"38", X"F1", --6D58
  X"CB", X"3F", X"30", X"0D", X"F5", X"EF", X"C1", X"E0", --6D60
  X"00", X"04", X"04", X"33", X"02", X"05", X"E1", X"38", --6D68
  X"F1", X"28", X"08", X"F5", X"EF", X"31", X"04", X"38", --6D70
  X"F1", X"18", X"E5", X"EF", X"02", X"38", X"C9", X"23", --6D78
  X"4E", X"23", X"7E", X"A9", X"91", X"5F", X"23", X"7E", --6D80
  X"89", X"A9", X"57", X"C9", X"0E", X"00", X"E5", X"36", --6D88
  X"00", X"23", X"71", X"23", X"7B", X"A9", X"91", X"77", --6D90
  X"23", X"7A", X"89", X"A9", X"77", X"23", X"36", X"00", --6D98
  X"E1", X"C9", X"EF", X"38", X"7E", X"A7", X"28", X"05", --6DA0
  X"EF", X"A2", X"0F", X"27", X"38", X"EF", X"02", X"38", --6DA8
  X"E5", X"D5", X"EB", X"46", X"CD", X"7F", X"2D", X"AF", --6DB0
  X"90", X"CB", X"79", X"42", X"4B", X"7B", X"D1", X"E1", --6DB8
  X"C9", X"57", X"17", X"9F", X"5F", X"4F", X"AF", X"47", --6DC0
  X"CD", X"B6", X"2A", X"EF", X"34", X"EF", X"1A", X"20", --6DC8
  X"9A", X"85", X"04", X"27", X"38", X"CD", X"A2", X"2D", --6DD0
  X"D8", X"F5", X"05", X"04", X"28", X"03", X"F1", X"37", --6DD8
  X"C9", X"F1", X"C9", X"EF", X"31", X"36", X"00", X"0B", --6DE0
  X"31", X"37", X"00", X"0D", X"02", X"38", X"3E", X"30", --6DE8
  X"D7", X"C9", X"2A", X"38", X"3E", X"2D", X"D7", X"EF", --6DF0
  X"A0", X"C3", X"C4", X"C5", X"02", X"38", X"D9", X"E5", --6DF8
  X"D9", X"EF", X"31", X"27", X"C2", X"03", X"E2", X"01", --6E00
  X"C2", X"02", X"38", X"7E", X"A7", X"20", X"47", X"CD", --6E08
  X"7F", X"2D", X"06", X"10", X"7A", X"A7", X"20", X"06", --6E10
  X"B3", X"28", X"09", X"53", X"06", X"08", X"D5", X"D9", --6E18
  X"D1", X"D9", X"18", X"57", X"EF", X"E2", X"38", X"7E", --6E20
  X"D6", X"7E", X"CD", X"C1", X"2D", X"57", X"3A", X"AC", --6E28
  X"5C", X"92", X"32", X"AC", X"5C", X"7A", X"CD", X"4F", --6E30
  X"2D", X"EF", X"31", X"27", X"C1", X"03", X"E1", X"38", --6E38
  X"CD", X"D5", X"2D", X"E5", X"32", X"A1", X"5C", X"3D", --6E40
  X"17", X"9F", X"3C", X"21", X"AB", X"5C", X"77", X"23", --6E48
  X"86", X"77", X"E1", X"C3", X"CF", X"2E", X"D6", X"80", --6E50
  X"FE", X"1C", X"38", X"13", X"CD", X"C1", X"2D", X"D6", --6E58
  X"07", X"47", X"21", X"AC", X"5C", X"86", X"77", X"78", --6E60
  X"ED", X"44", X"CD", X"4F", X"2D", X"18", X"92", X"EB", --6E68
  X"CD", X"BA", X"2F", X"D9", X"CB", X"FA", X"7D", X"D9", --6E70
  X"D6", X"80", X"47", X"CB", X"23", X"CB", X"12", X"D9", --6E78
  X"CB", X"13", X"CB", X"12", X"D9", X"21", X"AA", X"5C", --6E80
  X"0E", X"05", X"7E", X"8F", X"27", X"77", X"2B", X"0D", --6E88
  X"20", X"F8", X"10", X"E7", X"AF", X"21", X"A6", X"5C", --6E90
  X"11", X"A1", X"5C", X"06", X"09", X"ED", X"6F", X"0E", --6E98
  X"FF", X"ED", X"6F", X"20", X"04", X"0D", X"0C", X"20", --6EA0
  X"0A", X"12", X"13", X"FD", X"34", X"71", X"FD", X"34", --6EA8
  X"72", X"0E", X"00", X"CB", X"40", X"28", X"01", X"23", --6EB0
  X"10", X"E7", X"3A", X"AB", X"5C", X"D6", X"09", X"38", --6EB8
  X"0A", X"FD", X"35", X"71", X"3E", X"04", X"FD", X"BE", --6EC0
  X"6F", X"18", X"41", X"EF", X"02", X"E2", X"38", X"EB", --6EC8
  X"CD", X"BA", X"2F", X"D9", X"3E", X"80", X"95", X"2E", --6ED0
  X"00", X"CB", X"FA", X"D9", X"CD", X"DD", X"2F", X"FD", --6ED8
  X"7E", X"71", X"FE", X"08", X"38", X"06", X"D9", X"CB", --6EE0
  X"12", X"D9", X"18", X"20", X"01", X"00", X"02", X"7B", --6EE8
  X"CD", X"8B", X"2F", X"5F", X"7A", X"CD", X"8B", X"2F", --6EF0
  X"57", X"C5", X"D9", X"C1", X"10", X"F1", X"21", X"A1", --6EF8
  X"5C", X"79", X"FD", X"4E", X"71", X"09", X"77", X"FD", --6F00
  X"34", X"71", X"18", X"D3", X"F5", X"21", X"A1", X"5C", --6F08
  X"FD", X"4E", X"71", X"06", X"00", X"09", X"41", X"F1", --6F10
  X"2B", X"7E", X"CE", X"00", X"77", X"A7", X"28", X"05", --6F18
  X"FE", X"0A", X"3F", X"30", X"08", X"10", X"F1", X"36", --6F20
  X"01", X"04", X"FD", X"34", X"72", X"FD", X"70", X"71", --6F28
  X"EF", X"02", X"38", X"D9", X"E1", X"D9", X"ED", X"4B", --6F30
  X"AB", X"5C", X"21", X"A1", X"5C", X"78", X"FE", X"09", --6F38
  X"38", X"04", X"FE", X"FC", X"38", X"26", X"A7", X"CC", --6F40
  X"EF", X"15", X"AF", X"90", X"FA", X"52", X"2F", X"47", --6F48
  X"18", X"0C", X"79", X"A7", X"28", X"03", X"7E", X"23", --6F50
  X"0D", X"CD", X"EF", X"15", X"10", X"F4", X"79", X"A7", --6F58
  X"C8", X"04", X"3E", X"2E", X"D7", X"3E", X"30", X"10", --6F60
  X"FB", X"41", X"18", X"E6", X"50", X"15", X"06", X"01", --6F68
  X"CD", X"4A", X"2F", X"3E", X"45", X"D7", X"4A", X"79", --6F70
  X"A7", X"F2", X"83", X"2F", X"ED", X"44", X"4F", X"3E", --6F78
  X"2D", X"18", X"02", X"3E", X"2B", X"D7", X"06", X"00", --6F80
  X"C3", X"1B", X"1A", X"D5", X"6F", X"26", X"00", X"5D", --6F88
  X"54", X"29", X"29", X"19", X"29", X"59", X"19", X"4C", --6F90
  X"7D", X"D1", X"C9", X"7E", X"36", X"00", X"A7", X"C8", --6F98
  X"23", X"CB", X"7E", X"CB", X"FE", X"2B", X"C8", X"C5", --6FA0
  X"01", X"05", X"00", X"09", X"41", X"4F", X"37", X"2B", --6FA8
  X"7E", X"2F", X"CE", X"00", X"77", X"10", X"F8", X"79", --6FB0
  X"C1", X"C9", X"E5", X"F5", X"4E", X"23", X"46", X"77", --6FB8
  X"23", X"79", X"4E", X"C5", X"23", X"4E", X"23", X"46", --6FC0
  X"EB", X"57", X"5E", X"D5", X"23", X"56", X"23", X"5E", --6FC8
  X"D5", X"D9", X"D1", X"E1", X"C1", X"D9", X"23", X"56", --6FD0
  X"23", X"5E", X"F1", X"E1", X"C9", X"A7", X"C8", X"FE", --6FD8
  X"21", X"30", X"16", X"C5", X"47", X"D9", X"CB", X"2D", --6FE0
  X"CB", X"1A", X"CB", X"1B", X"D9", X"CB", X"1A", X"CB", --6FE8
  X"1B", X"10", X"F2", X"C1", X"D0", X"CD", X"04", X"30", --6FF0
  X"C0", X"D9", X"AF", X"2E", X"00", X"57", X"5D", X"D9", --6FF8
  X"11", X"00", X"00", X"C9", X"1C", X"C0", X"14", X"C0", --7000
  X"D9", X"1C", X"20", X"01", X"14", X"D9", X"C9", X"EB", --7008
  X"CD", X"6E", X"34", X"EB", X"1A", X"B6", X"20", X"26", --7010
  X"D5", X"23", X"E5", X"23", X"5E", X"23", X"56", X"23", --7018
  X"23", X"23", X"7E", X"23", X"4E", X"23", X"46", X"E1", --7020
  X"EB", X"09", X"EB", X"8E", X"0F", X"CE", X"00", X"20", --7028
  X"0B", X"9F", X"77", X"23", X"73", X"23", X"72", X"2B", --7030
  X"2B", X"2B", X"D1", X"C9", X"2B", X"D1", X"CD", X"93", --7038
  X"32", X"D9", X"E5", X"D9", X"D5", X"E5", X"CD", X"9B", --7040
  X"2F", X"47", X"EB", X"CD", X"9B", X"2F", X"4F", X"B8", --7048
  X"30", X"03", X"78", X"41", X"EB", X"F5", X"90", X"CD", --7050
  X"BA", X"2F", X"CD", X"DD", X"2F", X"F1", X"E1", X"77", --7058
  X"E5", X"68", X"61", X"19", X"D9", X"EB", X"ED", X"4A", --7060
  X"EB", X"7C", X"8D", X"6F", X"1F", X"AD", X"D9", X"EB", --7068
  X"E1", X"1F", X"30", X"08", X"3E", X"01", X"CD", X"DD", --7070
  X"2F", X"34", X"28", X"23", X"D9", X"7D", X"E6", X"80", --7078
  X"D9", X"23", X"77", X"2B", X"28", X"1F", X"7B", X"ED", --7080
  X"44", X"3F", X"5F", X"7A", X"2F", X"CE", X"00", X"57", --7088
  X"D9", X"7B", X"2F", X"CE", X"00", X"5F", X"7A", X"2F", --7090
  X"CE", X"00", X"30", X"07", X"1F", X"D9", X"34", X"CA", --7098
  X"AD", X"31", X"D9", X"57", X"D9", X"AF", X"C3", X"55", --70A0
  X"31", X"C5", X"06", X"10", X"7C", X"4D", X"21", X"00", --70A8
  X"00", X"29", X"38", X"0A", X"CB", X"11", X"17", X"30", --70B0
  X"03", X"19", X"38", X"02", X"10", X"F3", X"C1", X"C9", --70B8
  X"CD", X"E9", X"34", X"D8", X"23", X"AE", X"CB", X"FE", --70C0
  X"2B", X"C9", X"1A", X"B6", X"20", X"22", X"D5", X"E5", --70C8
  X"D5", X"CD", X"7F", X"2D", X"EB", X"E3", X"41", X"CD", --70D0
  X"7F", X"2D", X"78", X"A9", X"4F", X"E1", X"CD", X"A9", --70D8
  X"30", X"EB", X"E1", X"38", X"0A", X"7A", X"B3", X"20", --70E0
  X"01", X"4F", X"CD", X"8E", X"2D", X"D1", X"C9", X"D1", --70E8
  X"CD", X"93", X"32", X"AF", X"CD", X"C0", X"30", X"D8", --70F0
  X"D9", X"E5", X"D9", X"D5", X"EB", X"CD", X"C0", X"30", --70F8
  X"EB", X"38", X"5A", X"E5", X"CD", X"BA", X"2F", X"78", --7100
  X"A7", X"ED", X"62", X"D9", X"E5", X"ED", X"62", X"D9", --7108
  X"06", X"21", X"18", X"11", X"30", X"05", X"19", X"D9", --7110
  X"ED", X"5A", X"D9", X"D9", X"CB", X"1C", X"CB", X"1D", --7118
  X"D9", X"CB", X"1C", X"CB", X"1D", X"D9", X"CB", X"18", --7120
  X"CB", X"19", X"D9", X"CB", X"19", X"1F", X"10", X"E4", --7128
  X"EB", X"D9", X"EB", X"D9", X"C1", X"E1", X"78", X"81", --7130
  X"20", X"01", X"A7", X"3D", X"3F", X"17", X"3F", X"1F", --7138
  X"F2", X"46", X"31", X"30", X"68", X"A7", X"3C", X"20", --7140
  X"08", X"38", X"06", X"D9", X"CB", X"7A", X"D9", X"20", --7148
  X"5C", X"77", X"D9", X"78", X"D9", X"30", X"15", X"7E", --7150
  X"A7", X"3E", X"80", X"28", X"01", X"AF", X"D9", X"A2", --7158
  X"CD", X"FB", X"2F", X"07", X"77", X"38", X"2E", X"23", --7160
  X"77", X"2B", X"18", X"29", X"06", X"20", X"D9", X"CB", --7168
  X"7A", X"D9", X"20", X"12", X"07", X"CB", X"13", X"CB", --7170
  X"12", X"D9", X"CB", X"13", X"CB", X"12", X"D9", X"35", --7178
  X"28", X"D7", X"10", X"EA", X"18", X"D7", X"17", X"30", --7180
  X"0C", X"CD", X"04", X"30", X"20", X"07", X"D9", X"16", --7188
  X"80", X"D9", X"34", X"28", X"18", X"E5", X"23", X"D9", --7190
  X"D5", X"D9", X"C1", X"78", X"17", X"CB", X"16", X"1F", --7198
  X"77", X"23", X"71", X"23", X"72", X"23", X"73", X"E1", --71A0
  X"D1", X"D9", X"E1", X"D9", X"C9", X"CF", X"05", X"CD", --71A8
  X"93", X"32", X"EB", X"AF", X"CD", X"C0", X"30", X"38", --71B0
  X"F4", X"EB", X"CD", X"C0", X"30", X"D8", X"D9", X"E5", --71B8
  X"D9", X"D5", X"E5", X"CD", X"BA", X"2F", X"D9", X"E5", --71C0
  X"60", X"69", X"D9", X"61", X"68", X"AF", X"06", X"DF", --71C8
  X"18", X"10", X"17", X"CB", X"11", X"D9", X"CB", X"11", --71D0
  X"CB", X"10", X"D9", X"29", X"D9", X"ED", X"6A", X"D9", --71D8
  X"38", X"10", X"ED", X"52", X"D9", X"ED", X"52", X"D9", --71E0
  X"30", X"0F", X"19", X"D9", X"ED", X"5A", X"D9", X"A7", --71E8
  X"18", X"08", X"A7", X"ED", X"52", X"D9", X"ED", X"52", --71F0
  X"D9", X"37", X"04", X"FA", X"D2", X"31", X"F5", X"28", --71F8
  X"E1", X"5F", X"51", X"D9", X"59", X"50", X"F1", X"CB", --7200
  X"18", X"F1", X"CB", X"18", X"D9", X"C1", X"E1", X"78", --7208
  X"91", X"C3", X"3D", X"31", X"7E", X"A7", X"C8", X"FE", --7210
  X"81", X"30", X"06", X"36", X"00", X"3E", X"20", X"18", --7218
  X"51", X"FE", X"91", X"20", X"1A", X"23", X"23", X"23", --7220
  X"3E", X"80", X"A6", X"2B", X"B6", X"2B", X"20", X"03", --7228
  X"3E", X"80", X"AE", X"2B", X"20", X"36", X"77", X"23", --7230
  X"36", X"FF", X"2B", X"3E", X"18", X"18", X"33", X"30", --7238
  X"2C", X"D5", X"2F", X"C6", X"91", X"23", X"56", X"23", --7240
  X"5E", X"2B", X"2B", X"0E", X"00", X"CB", X"7A", X"28", --7248
  X"01", X"0D", X"CB", X"FA", X"06", X"08", X"90", X"80", --7250
  X"38", X"04", X"5A", X"16", X"00", X"90", X"28", X"07", --7258
  X"47", X"CB", X"3A", X"CB", X"1B", X"10", X"FA", X"CD", --7260
  X"8E", X"2D", X"D1", X"C9", X"7E", X"D6", X"A0", X"F0", --7268
  X"ED", X"44", X"D5", X"EB", X"2B", X"47", X"CB", X"38", --7270
  X"CB", X"38", X"CB", X"38", X"28", X"05", X"36", X"00", --7278
  X"2B", X"10", X"FB", X"E6", X"07", X"28", X"09", X"47", --7280
  X"3E", X"FF", X"CB", X"27", X"10", X"FC", X"A6", X"77", --7288
  X"EB", X"D1", X"C9", X"CD", X"96", X"32", X"EB", X"7E", --7290
  X"A7", X"C0", X"D5", X"CD", X"7F", X"2D", X"AF", X"23", --7298
  X"77", X"2B", X"77", X"06", X"91", X"7A", X"A7", X"20", --72A0
  X"08", X"B3", X"42", X"28", X"10", X"53", X"58", X"06", --72A8
  X"89", X"EB", X"05", X"29", X"30", X"FC", X"CB", X"09", --72B0
  X"CB", X"1C", X"CB", X"1D", X"EB", X"2B", X"73", X"2B", --72B8
  X"72", X"2B", X"70", X"D1", X"C9", X"00", X"B0", X"00", --72C0
  X"40", X"B0", X"00", X"01", X"30", X"00", X"F1", X"49", --72C8
  X"0F", X"DA", X"A2", X"40", X"B0", X"00", X"0A", X"8F", --72D0
  X"36", X"3C", X"34", X"A1", X"33", X"0F", X"30", X"CA", --72D8
  X"30", X"AF", X"31", X"51", X"38", X"1B", X"35", X"24", --72E0
  X"35", X"3B", X"35", X"3B", X"35", X"3B", X"35", X"3B", --72E8
  X"35", X"3B", X"35", X"3B", X"35", X"14", X"30", X"2D", --72F0
  X"35", X"3B", X"35", X"3B", X"35", X"3B", X"35", X"3B", --72F8
  X"35", X"3B", X"35", X"3B", X"35", X"9C", X"35", X"DE", --7300
  X"35", X"BC", X"34", X"45", X"36", X"6E", X"34", X"69", --7308
  X"36", X"DE", X"35", X"74", X"36", X"B5", X"37", X"AA", --7310
  X"37", X"DA", X"37", X"33", X"38", X"43", X"38", X"E2", --7318
  X"37", X"13", X"37", X"C4", X"36", X"AF", X"36", X"4A", --7320
  X"38", X"92", X"34", X"6A", X"34", X"AC", X"34", X"A5", --7328
  X"34", X"B3", X"34", X"1F", X"36", X"C9", X"35", X"01", --7330
  X"35", X"C0", X"33", X"A0", X"36", X"86", X"36", X"C6", --7338
  X"33", X"7A", X"36", X"06", X"35", X"F9", X"34", X"9B", --7340
  X"36", X"83", X"37", X"14", X"32", X"A2", X"33", X"4F", --7348
  X"2D", X"97", X"32", X"49", X"34", X"1B", X"34", X"2D", --7350
  X"34", X"0F", X"34", X"CD", X"BF", X"35", X"78", X"32", --7358
  X"67", X"5C", X"D9", X"E3", X"D9", X"ED", X"53", X"65", --7360
  X"5C", X"D9", X"7E", X"23", X"E5", X"A7", X"F2", X"80", --7368
  X"33", X"57", X"E6", X"60", X"0F", X"0F", X"0F", X"0F", --7370
  X"C6", X"7C", X"6F", X"7A", X"E6", X"1F", X"18", X"0E", --7378
  X"FE", X"18", X"30", X"08", X"D9", X"01", X"FB", X"FF", --7380
  X"54", X"5D", X"09", X"D9", X"07", X"6F", X"11", X"D7", --7388
  X"32", X"26", X"00", X"19", X"5E", X"23", X"56", X"21", --7390
  X"65", X"33", X"E3", X"D5", X"D9", X"ED", X"4B", X"66", --7398
  X"5C", X"C9", X"F1", X"3A", X"67", X"5C", X"D9", X"18", --73A0
  X"C3", X"D5", X"E5", X"01", X"05", X"00", X"CD", X"05", --73A8
  X"1F", X"E1", X"D1", X"C9", X"ED", X"5B", X"65", X"5C", --73B0
  X"CD", X"C0", X"33", X"ED", X"53", X"65", X"5C", X"C9", --73B8
  X"CD", X"A9", X"33", X"ED", X"B0", X"C9", X"62", X"6B", --73C0
  X"CD", X"A9", X"33", X"D9", X"E5", X"D9", X"E3", X"C5", --73C8
  X"7E", X"E6", X"C0", X"07", X"07", X"4F", X"0C", X"7E", --73D0
  X"E6", X"3F", X"20", X"02", X"23", X"7E", X"C6", X"50", --73D8
  X"12", X"3E", X"05", X"91", X"23", X"13", X"06", X"00", --73E0
  X"ED", X"B0", X"C1", X"E3", X"D9", X"E1", X"D9", X"47", --73E8
  X"AF", X"05", X"C8", X"12", X"13", X"18", X"FA", X"A7", --73F0
  X"C8", X"F5", X"D5", X"11", X"00", X"00", X"CD", X"C8", --73F8
  X"33", X"D1", X"F1", X"3D", X"18", X"F2", X"4F", X"07", --7400
  X"07", X"81", X"4F", X"06", X"00", X"09", X"C9", X"D5", --7408
  X"2A", X"68", X"5C", X"CD", X"06", X"34", X"CD", X"C0", --7410
  X"33", X"E1", X"C9", X"62", X"6B", X"D9", X"E5", X"21", --7418
  X"C5", X"32", X"D9", X"CD", X"F7", X"33", X"CD", X"C8", --7420
  X"33", X"D9", X"E1", X"D9", X"C9", X"E5", X"EB", X"2A", --7428
  X"68", X"5C", X"CD", X"06", X"34", X"EB", X"CD", X"C0", --7430
  X"33", X"EB", X"E1", X"C9", X"06", X"05", X"1A", X"4E", --7438
  X"EB", X"12", X"71", X"23", X"13", X"10", X"F7", X"EB", --7440
  X"C9", X"47", X"CD", X"5E", X"33", X"31", X"0F", X"C0", --7448
  X"02", X"A0", X"C2", X"31", X"E0", X"04", X"E2", X"C1", --7450
  X"03", X"38", X"CD", X"C6", X"33", X"CD", X"62", X"33", --7458
  X"0F", X"01", X"C2", X"02", X"35", X"EE", X"E1", X"03", --7460
  X"38", X"C9", X"06", X"FF", X"18", X"06", X"CD", X"E9", --7468
  X"34", X"D8", X"06", X"00", X"7E", X"A7", X"28", X"0B", --7470
  X"23", X"78", X"E6", X"80", X"B6", X"17", X"3F", X"1F", --7478
  X"77", X"2B", X"C9", X"D5", X"E5", X"CD", X"7F", X"2D", --7480
  X"E1", X"78", X"B1", X"2F", X"4F", X"CD", X"8E", X"2D", --7488
  X"D1", X"C9", X"CD", X"E9", X"34", X"D8", X"D5", X"11", --7490
  X"01", X"00", X"23", X"CB", X"16", X"2B", X"9F", X"4F", --7498
  X"CD", X"8E", X"2D", X"D1", X"C9", X"CD", X"99", X"1E", --74A0
  X"ED", X"78", X"18", X"04", X"CD", X"99", X"1E", X"0A", --74A8
  X"C3", X"28", X"2D", X"CD", X"99", X"1E", X"21", X"2B", --74B0
  X"2D", X"E5", X"C5", X"C9", X"CD", X"F1", X"2B", X"0B", --74B8
  X"78", X"B1", X"20", X"23", X"1A", X"CD", X"8D", X"2C", --74C0
  X"38", X"09", X"D6", X"90", X"38", X"19", X"FE", X"15", --74C8
  X"30", X"15", X"3C", X"3D", X"87", X"87", X"87", X"FE", --74D0
  X"A8", X"30", X"0C", X"ED", X"4B", X"7B", X"5C", X"81", --74D8
  X"4F", X"30", X"01", X"04", X"C3", X"2B", X"2D", X"CF", --74E0
  X"09", X"E5", X"C5", X"47", X"7E", X"23", X"B6", X"23", --74E8
  X"B6", X"23", X"B6", X"78", X"C1", X"E1", X"C0", X"37", --74F0
  X"C9", X"CD", X"E9", X"34", X"D8", X"3E", X"FF", X"18", --74F8
  X"06", X"CD", X"E9", X"34", X"18", X"05", X"AF", X"23", --7500
  X"AE", X"2B", X"07", X"E5", X"3E", X"00", X"77", X"23", --7508
  X"77", X"23", X"17", X"77", X"1F", X"23", X"77", X"23", --7510
  X"77", X"E1", X"C9", X"EB", X"CD", X"E9", X"34", X"EB", --7518
  X"D8", X"37", X"18", X"E7", X"EB", X"CD", X"E9", X"34", --7520
  X"EB", X"D0", X"A7", X"18", X"DE", X"EB", X"CD", X"E9", --7528
  X"34", X"EB", X"D0", X"D5", X"1B", X"AF", X"12", X"1B", --7530
  X"12", X"D1", X"C9", X"78", X"D6", X"08", X"CB", X"57", --7538
  X"20", X"01", X"3D", X"0F", X"30", X"08", X"F5", X"E5", --7540
  X"CD", X"3C", X"34", X"D1", X"EB", X"F1", X"CB", X"57", --7548
  X"20", X"07", X"0F", X"F5", X"CD", X"0F", X"30", X"18", --7550
  X"33", X"0F", X"F5", X"CD", X"F1", X"2B", X"D5", X"C5", --7558
  X"CD", X"F1", X"2B", X"E1", X"7C", X"B5", X"E3", X"78", --7560
  X"20", X"0B", X"B1", X"C1", X"28", X"04", X"F1", X"3F", --7568
  X"18", X"16", X"F1", X"18", X"13", X"B1", X"28", X"0D", --7570
  X"1A", X"96", X"38", X"09", X"20", X"ED", X"0B", X"13", --7578
  X"23", X"E3", X"2B", X"18", X"DF", X"C1", X"F1", X"A7", --7580
  X"F5", X"EF", X"A0", X"38", X"F1", X"F5", X"DC", X"01", --7588
  X"35", X"F1", X"F5", X"D4", X"F9", X"34", X"F1", X"0F", --7590
  X"D4", X"01", X"35", X"C9", X"CD", X"F1", X"2B", X"D5", --7598
  X"C5", X"CD", X"F1", X"2B", X"E1", X"E5", X"D5", X"C5", --75A0
  X"09", X"44", X"4D", X"F7", X"CD", X"B2", X"2A", X"C1", --75A8
  X"E1", X"78", X"B1", X"28", X"02", X"ED", X"B0", X"C1", --75B0
  X"E1", X"78", X"B1", X"28", X"02", X"ED", X"B0", X"2A", --75B8
  X"65", X"5C", X"11", X"FB", X"FF", X"E5", X"19", X"D1", --75C0
  X"C9", X"CD", X"D5", X"2D", X"38", X"0E", X"20", X"0C", --75C8
  X"F5", X"01", X"01", X"00", X"F7", X"F1", X"12", X"CD", --75D0
  X"B2", X"2A", X"EB", X"C9", X"CF", X"0A", X"2A", X"5D", --75D8
  X"5C", X"E5", X"78", X"C6", X"E3", X"9F", X"F5", X"CD", --75E0
  X"F1", X"2B", X"D5", X"03", X"F7", X"E1", X"ED", X"53", --75E8
  X"5D", X"5C", X"D5", X"ED", X"B0", X"EB", X"2B", X"36", --75F0
  X"0D", X"FD", X"CB", X"01", X"BE", X"CD", X"FB", X"24", --75F8
  X"DF", X"FE", X"0D", X"20", X"07", X"E1", X"F1", X"FD", --7600
  X"AE", X"01", X"E6", X"40", X"C2", X"8A", X"1C", X"22", --7608
  X"5D", X"5C", X"FD", X"CB", X"01", X"FE", X"CD", X"FB", --7610
  X"24", X"E1", X"22", X"5D", X"5C", X"18", X"A0", X"01", --7618
  X"01", X"00", X"F7", X"22", X"5B", X"5C", X"E5", X"2A", --7620
  X"51", X"5C", X"E5", X"3E", X"FF", X"CD", X"01", X"16", --7628
  X"CD", X"E3", X"2D", X"E1", X"CD", X"15", X"16", X"D1", --7630
  X"2A", X"5B", X"5C", X"A7", X"ED", X"52", X"44", X"4D", --7638
  X"CD", X"B2", X"2A", X"EB", X"C9", X"CD", X"94", X"1E", --7640
  X"FE", X"10", X"D2", X"9F", X"1E", X"2A", X"51", X"5C", --7648
  X"E5", X"CD", X"01", X"16", X"CD", X"E6", X"15", X"01", --7650
  X"00", X"00", X"30", X"03", X"0C", X"F7", X"12", X"CD", --7658
  X"B2", X"2A", X"E1", X"CD", X"15", X"16", X"C3", X"BF", --7660
  X"35", X"CD", X"F1", X"2B", X"78", X"B1", X"28", X"01", --7668
  X"1A", X"C3", X"28", X"2D", X"CD", X"F1", X"2B", X"C3", --7670
  X"2B", X"2D", X"D9", X"E5", X"21", X"67", X"5C", X"35", --7678
  X"E1", X"20", X"04", X"23", X"D9", X"C9", X"D9", X"5E", --7680
  X"7B", X"17", X"9F", X"57", X"19", X"D9", X"C9", X"13", --7688
  X"13", X"1A", X"1B", X"1B", X"A7", X"20", X"EF", X"D9", --7690
  X"23", X"D9", X"C9", X"F1", X"D9", X"E3", X"D9", X"C9", --7698
  X"EF", X"C0", X"02", X"31", X"E0", X"05", X"27", X"E0", --76A0
  X"01", X"C0", X"04", X"03", X"E0", X"38", X"C9", X"EF", --76A8
  X"31", X"36", X"00", X"04", X"3A", X"38", X"C9", X"31", --76B0
  X"3A", X"C0", X"03", X"E0", X"01", X"30", X"00", X"03", --76B8
  X"A1", X"03", X"38", X"C9", X"EF", X"3D", X"34", X"F1", --76C0
  X"38", X"AA", X"3B", X"29", X"04", X"31", X"27", X"C3", --76C8
  X"03", X"31", X"0F", X"A1", X"03", X"88", X"13", X"36", --76D0
  X"58", X"65", X"66", X"9D", X"78", X"65", X"40", X"A2", --76D8
  X"60", X"32", X"C9", X"E7", X"21", X"F7", X"AF", X"24", --76E0
  X"EB", X"2F", X"B0", X"B0", X"14", X"EE", X"7E", X"BB", --76E8
  X"94", X"58", X"F1", X"3A", X"7E", X"F8", X"CF", X"E3", --76F0
  X"38", X"CD", X"D5", X"2D", X"20", X"07", X"38", X"03", --76F8
  X"86", X"30", X"09", X"CF", X"05", X"38", X"07", X"96", --7700
  X"30", X"04", X"ED", X"44", X"77", X"C9", X"EF", X"02", --7708
  X"A0", X"38", X"C9", X"EF", X"3D", X"31", X"37", X"00", --7710
  X"04", X"38", X"CF", X"09", X"A0", X"02", X"38", X"7E", --7718
  X"36", X"80", X"CD", X"28", X"2D", X"EF", X"34", X"38", --7720
  X"00", X"03", X"01", X"31", X"34", X"F0", X"4C", X"CC", --7728
  X"CC", X"CD", X"03", X"37", X"00", X"08", X"01", X"A1", --7730
  X"03", X"01", X"38", X"34", X"EF", X"01", X"34", X"F0", --7738
  X"31", X"72", X"17", X"F8", X"04", X"01", X"A2", X"03", --7740
  X"A2", X"03", X"31", X"34", X"32", X"20", X"04", X"A2", --7748
  X"03", X"8C", X"11", X"AC", X"14", X"09", X"56", X"DA", --7750
  X"A5", X"59", X"30", X"C5", X"5C", X"90", X"AA", X"9E", --7758
  X"70", X"6F", X"61", X"A1", X"CB", X"DA", X"96", X"A4", --7760
  X"31", X"9F", X"B4", X"E7", X"A0", X"FE", X"5C", X"FC", --7768
  X"EA", X"1B", X"43", X"CA", X"36", X"ED", X"A7", X"9C", --7770
  X"7E", X"5E", X"F0", X"6E", X"23", X"80", X"93", X"04", --7778
  X"0F", X"38", X"C9", X"EF", X"3D", X"34", X"EE", X"22", --7780
  X"F9", X"83", X"6E", X"04", X"31", X"A2", X"0F", X"27", --7788
  X"03", X"31", X"0F", X"31", X"0F", X"31", X"2A", X"A1", --7790
  X"03", X"31", X"37", X"C0", X"00", X"04", X"02", X"38", --7798
  X"C9", X"A1", X"03", X"01", X"36", X"00", X"02", X"1B", --77A0
  X"38", X"C9", X"EF", X"39", X"2A", X"A1", X"03", X"E0", --77A8
  X"00", X"06", X"1B", X"33", X"03", X"EF", X"39", X"31", --77B0
  X"31", X"04", X"31", X"0F", X"A1", X"03", X"86", X"14", --77B8
  X"E6", X"5C", X"1F", X"0B", X"A3", X"8F", X"38", X"EE", --77C0
  X"E9", X"15", X"63", X"BB", X"23", X"EE", X"92", X"0D", --77C8
  X"CD", X"ED", X"F1", X"23", X"5D", X"1B", X"EA", X"04", --77D0
  X"38", X"C9", X"EF", X"31", X"1F", X"01", X"20", X"05", --77D8
  X"38", X"C9", X"CD", X"97", X"32", X"7E", X"FE", X"81", --77E0
  X"38", X"0E", X"EF", X"A1", X"1B", X"01", X"05", X"31", --77E8
  X"36", X"A3", X"01", X"00", X"06", X"1B", X"33", X"03", --77F0
  X"EF", X"A0", X"01", X"31", X"31", X"04", X"31", X"0F", --77F8
  X"A1", X"03", X"8C", X"10", X"B2", X"13", X"0E", X"55", --7800
  X"E4", X"8D", X"58", X"39", X"BC", X"5B", X"98", X"FD", --7808
  X"9E", X"00", X"36", X"75", X"A0", X"DB", X"E8", X"B4", --7810
  X"63", X"42", X"C4", X"E6", X"B5", X"09", X"36", X"BE", --7818
  X"E9", X"36", X"73", X"1B", X"5D", X"EC", X"D8", X"DE", --7820
  X"63", X"BE", X"F0", X"61", X"A1", X"B3", X"0C", X"04", --7828
  X"0F", X"38", X"C9", X"EF", X"31", X"31", X"04", X"A1", --7830
  X"03", X"1B", X"28", X"A1", X"0F", X"05", X"24", X"31", --7838
  X"0F", X"38", X"C9", X"EF", X"22", X"A3", X"03", X"1B", --7840
  X"38", X"C9", X"EF", X"31", X"30", X"00", X"1E", X"A2", --7848
  X"38", X"EF", X"01", X"31", X"30", X"00", X"07", X"25", --7850
  X"04", X"38", X"C3", X"C4", X"36", X"02", X"31", X"30", --7858
  X"00", X"09", X"A0", X"01", X"37", X"00", X"06", X"A1", --7860
  X"01", X"05", X"02", X"A1", X"38", X"C9", X"DD", X"E5", --7868
  X"FD", X"CB", X"01", X"66", X"28", X"03", X"CD", X"42", --7870
  X"3A", X"CD", X"BF", X"02", X"DD", X"E1", X"C9", X"0E", --7878
  X"FD", X"16", X"FF", X"1E", X"BF", X"42", X"3E", X"07", --7880
  X"ED", X"79", X"ED", X"60", X"3E", X"0E", X"ED", X"79", --7888
  X"ED", X"78", X"F6", X"F0", X"6F", X"C9", X"42", X"3E", --7890
  X"0E", X"ED", X"79", X"43", X"ED", X"69", X"C9", X"42", --7898
  X"3E", X"0E", X"ED", X"79", X"ED", X"78", X"C9", X"7D", --78A0
  X"E6", X"FE", X"6F", X"18", X"E9", X"7D", X"F6", X"01", --78A8
  X"6F", X"18", X"E3", X"10", X"FE", X"C9", X"C5", X"06", --78B0
  X"10", X"CD", X"B3", X"38", X"C1", X"10", X"F7", X"C9", --78B8
  X"C5", X"CD", X"9F", X"38", X"C1", X"E6", X"20", X"28", --78C0
  X"02", X"10", X"F5", X"C9", X"C5", X"CD", X"9F", X"38", --78C8
  X"C1", X"E6", X"20", X"20", X"02", X"10", X"F5", X"C9", --78D0
  X"CD", X"7F", X"38", X"06", X"01", X"18", X"05", X"CD", --78D8
  X"7F", X"38", X"06", X"04", X"C5", X"CD", X"9F", X"38", --78E0
  X"C1", X"E6", X"20", X"28", X"40", X"AF", X"C5", X"F5", --78E8
  X"CD", X"AD", X"38", X"06", X"A3", X"CD", X"C0", X"38", --78F0
  X"20", X"31", X"CD", X"A7", X"38", X"18", X"02", X"FF", --78F8
  X"FF", X"06", X"2B", X"CD", X"B3", X"38", X"CD", X"9F", --7900
  X"38", X"CB", X"6F", X"28", X"04", X"F1", X"37", X"18", --7908
  X"03", X"F1", X"37", X"3F", X"1F", X"F5", X"CD", X"AD", --7910
  X"38", X"06", X"26", X"CD", X"B3", X"38", X"CD", X"A7", --7918
  X"38", X"06", X"23", X"CD", X"B3", X"38", X"F1", X"C1", --7920
  X"10", X"C4", X"C9", X"F1", X"C1", X"CD", X"AD", X"38", --7928
  X"AF", X"32", X"88", X"5B", X"3C", X"37", X"3F", X"C9", --7930
  X"CD", X"7F", X"38", X"3A", X"88", X"5B", X"E6", X"80", --7938
  X"20", X"57", X"CD", X"9F", X"38", X"E6", X"20", X"28", --7940
  X"E4", X"3A", X"88", X"5B", X"A7", X"20", X"0B", X"3C", --7948
  X"32", X"88", X"5B", X"3E", X"4C", X"32", X"89", X"5B", --7950
  X"18", X"42", X"3A", X"89", X"5B", X"3D", X"32", X"89", --7958
  X"5B", X"20", X"39", X"AF", X"32", X"88", X"5B", X"32", --7960
  X"89", X"5B", X"32", X"8A", X"5B", X"CD", X"A7", X"38", --7968
  X"06", X"21", X"CD", X"C0", X"38", X"20", X"B6", X"CD", --7970
  X"AD", X"38", X"06", X"24", X"CD", X"CC", X"38", X"28", --7978
  X"AC", X"CD", X"A7", X"38", X"06", X"0F", X"CD", X"B6", --7980
  X"38", X"CD", X"DF", X"38", X"20", X"9F", X"CB", X"FF", --7988
  X"E6", X"F0", X"32", X"88", X"5B", X"AF", X"CB", X"3F", --7990
  X"C9", X"AF", X"37", X"C9", X"AF", X"3C", X"37", X"C9", --7998
  X"CD", X"38", X"39", X"3A", X"88", X"5B", X"2F", X"E6", --79A0
  X"C0", X"C0", X"DD", X"21", X"8A", X"5B", X"06", X"05", --79A8
  X"C5", X"CD", X"D8", X"38", X"C2", X"3A", X"3A", X"CB", --79B0
  X"7F", X"28", X"21", X"CD", X"DF", X"38", X"20", X"7A", --79B8
  X"C1", X"C5", X"4F", X"DD", X"7E", X"00", X"CB", X"40", --79C0
  X"28", X"0C", X"CB", X"39", X"CB", X"39", X"CB", X"39", --79C8
  X"CB", X"39", X"E6", X"F0", X"18", X"02", X"E6", X"0F", --79D0
  X"B1", X"DD", X"77", X"00", X"C1", X"CB", X"40", X"20", --79D8
  X"02", X"DD", X"2B", X"10", X"CB", X"1E", X"80", X"DD", --79E0
  X"21", X"88", X"5B", X"21", X"3F", X"3A", X"06", X"03", --79E8
  X"DD", X"7E", X"00", X"A6", X"28", X"21", X"CB", X"7B", --79F0
  X"28", X"42", X"C5", X"F5", X"78", X"18", X"02", X"FF", --79F8
  X"FF", X"3D", X"CB", X"27", X"CB", X"27", X"CB", X"27", --7A00
  X"F6", X"07", X"47", X"F1", X"CB", X"27", X"DA", X"13", --7A08
  X"3A", X"10", X"F9", X"58", X"C1", X"20", X"25", X"DD", --7A10
  X"23", X"23", X"10", X"D4", X"CB", X"7B", X"20", X"07", --7A18
  X"7B", X"E6", X"FC", X"28", X"02", X"1D", X"1D", X"3A", --7A20
  X"8A", X"5B", X"E6", X"08", X"28", X"06", X"7B", X"E6", --7A28
  X"7F", X"C6", X"12", X"5F", X"7B", X"C6", X"5A", X"5F", --7A30
  X"AF", X"C9", X"C1", X"C9", X"AF", X"3C", X"C9", X"0F", --7A38
  X"FF", X"F2", X"1E", X"80", X"3A", X"78", X"5C", X"E6", --7A40
  X"01", X"20", X"04", X"CD", X"A0", X"39", X"C0", X"21", --7A48
  X"00", X"5C", X"CB", X"7E", X"20", X"0C", X"7E", X"FE", --7A50
  X"5B", X"38", X"07", X"23", X"35", X"2B", X"20", X"02", --7A58
  X"36", X"FF", X"7D", X"21", X"04", X"5C", X"BD", X"20", --7A60
  X"E9", X"CD", X"AE", X"3A", X"C0", X"7B", X"21", X"00", --7A68
  X"5C", X"BE", X"28", X"2A", X"EB", X"21", X"04", X"5C", --7A70
  X"BE", X"28", X"23", X"CB", X"7E", X"20", X"04", X"EB", --7A78
  X"CB", X"7E", X"C8", X"5F", X"77", X"23", X"36", X"0A", --7A80
  X"23", X"3A", X"09", X"5C", X"CB", X"3F", X"77", X"23", --7A88
  X"CD", X"D7", X"3A", X"73", X"7B", X"32", X"08", X"5C", --7A90
  X"21", X"3B", X"5C", X"CB", X"EE", X"C9", X"23", X"36", --7A98
  X"0A", X"23", X"35", X"C0", X"3A", X"0A", X"5C", X"CB", --7AA0
  X"3F", X"77", X"23", X"5E", X"18", X"E6", X"7B", X"21", --7AA8
  X"66", X"5B", X"CB", X"46", X"28", X"06", X"FE", X"6D", --7AB0
  X"30", X"1A", X"AF", X"C9", X"FE", X"80", X"30", X"14", --7AB8
  X"FE", X"6C", X"20", X"F6", X"00", X"00", X"00", X"00", --7AC0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --7AC8
  X"00", X"00", X"00", X"00", X"AF", X"3C", X"C9", X"E5", --7AD0
  X"7B", X"D6", X"5B", X"16", X"00", X"5F", X"21", X"66", --7AD8
  X"5B", X"CB", X"46", X"28", X"05", X"21", X"13", X"3B", --7AE0
  X"18", X"25", X"21", X"25", X"3B", X"FE", X"11", X"38", --7AE8
  X"1E", X"21", X"21", X"3B", X"FE", X"15", X"28", X"17", --7AF0
  X"FE", X"16", X"28", X"13", X"18", X"03", X"00", X"FF", --7AF8
  X"FF", X"FE", X"17", X"28", X"0A", X"21", X"18", X"3B", --7B00
  X"FE", X"21", X"30", X"03", X"21", X"13", X"3B", X"19", --7B08
  X"5E", X"E1", X"C9", X"2E", X"0D", X"33", X"32", X"31", --7B10
  X"29", X"28", X"2A", X"2F", X"2D", X"39", X"38", X"37", --7B18
  X"2B", X"36", X"35", X"34", X"30", X"A5", X"0D", X"A6", --7B20
  X"A7", X"A8", X"A9", X"AA", X"0B", X"0C", X"07", X"09", --7B28
  X"0A", X"08", X"AC", X"AD", X"AE", X"AF", X"B0", X"B1", --7B30
  X"B2", X"B3", X"B4", X"FD", X"CB", X"01", X"66", X"20", --7B38
  X"05", X"AF", X"11", X"36", X"15", X"C9", X"21", X"0F", --7B40
  X"01", X"E3", X"C3", X"00", X"5B", X"FD", X"CB", X"01", --7B48
  X"66", X"20", X"05", X"FD", X"CB", X"0A", X"7E", X"C9", --7B50
  X"21", X"12", X"01", X"18", X"EC", X"FD", X"CB", X"01", --7B58
  X"66", X"20", X"04", X"DF", X"FE", X"0D", X"C9", X"21", --7B60
  X"15", X"01", X"18", X"DD", X"CD", X"8E", X"02", X"0E", --7B68
  X"00", X"20", X"0D", X"CD", X"1E", X"03", X"30", X"08", --7B70
  X"15", X"5F", X"CD", X"33", X"03", X"C3", X"57", X"26", --7B78
  X"FD", X"CB", X"01", X"66", X"CA", X"60", X"26", X"F3", --7B80
  X"CD", X"A0", X"39", X"FB", X"20", X"0C", X"CD", X"AE", --7B88
  X"3A", X"20", X"07", X"CD", X"D7", X"3A", X"7B", X"C3", --7B90
  X"57", X"26", X"0E", X"00", X"C3", X"60", X"26", X"FE", --7B98
  X"A3", X"28", X"0C", X"FE", X"A4", X"28", X"08", X"D6", --7BA0
  X"A5", X"D2", X"5F", X"0B", X"C3", X"56", X"0B", X"FD", --7BA8
  X"CB", X"01", X"66", X"28", X"F2", X"11", X"C9", X"3B", --7BB0
  X"D5", X"D6", X"A3", X"11", X"D2", X"3B", X"28", X"03", --7BB8
  X"11", X"DA", X"3B", X"3E", X"04", X"F5", X"C3", X"17", --7BC0
  X"0C", X"37", X"FD", X"CB", X"01", X"4E", X"C0", X"C3", --7BC8
  X"03", X"0B", X"53", X"50", X"45", X"43", X"54", X"52", --7BD0
  X"55", X"CD", X"50", X"4C", X"41", X"D9", X"C3", X"01", --7BD8
  X"3C", X"69", X"51", X"59", X"ED", X"B0", X"01", X"FD", --7BE0
  X"7F", X"3E", X"07", X"ED", X"79", X"26", X"C0", X"54", --7BE8
  X"01", X"00", X"40", X"ED", X"B0", X"1B", X"AF", X"01", --7BF0
  X"FD", X"7F", X"ED", X"79", X"C3", X"CB", X"11", X"FF", --7BF8
  X"FF", X"C3", X"A0", X"39", X"C3", X"10", X"3C", X"C3", --7C00
  X"10", X"3C", X"C3", X"10", X"3C", X"C3", X"10", X"3C", --7C08
  X"3E", X"7F", X"DB", X"FE", X"1F", X"D8", X"3E", X"FE", --7C10
  X"DB", X"FE", X"1F", X"D8", X"3E", X"07", X"D3", X"FE", --7C18
  X"3E", X"02", X"CD", X"01", X"16", X"AF", X"32", X"3C", --7C20
  X"5C", X"3E", X"16", X"D7", X"AF", X"D7", X"AF", X"D7", --7C28
  X"1E", X"08", X"43", X"50", X"78", X"3D", X"CB", X"17", --7C30
  X"CB", X"17", X"CB", X"17", X"82", X"3D", X"32", X"8F", --7C38
  X"5C", X"21", X"8F", X"3C", X"4B", X"7E", X"D7", X"23", --7C40
  X"0D", X"20", X"FA", X"10", X"E7", X"43", X"15", X"20", --7C48
  X"E3", X"21", X"00", X"48", X"54", X"5D", X"13", X"AF", --7C50
  X"77", X"01", X"FF", X"0F", X"ED", X"B0", X"EB", X"11", --7C58
  X"00", X"59", X"01", X"00", X"02", X"ED", X"B0", X"F3", --7C60
  X"11", X"70", X"03", X"2E", X"07", X"01", X"99", X"00", --7C68
  X"0B", X"78", X"B1", X"20", X"FB", X"7D", X"EE", X"10", --7C70
  X"6F", X"D3", X"FE", X"1B", X"7A", X"B3", X"20", X"ED", --7C78
  X"01", X"00", X"00", X"0B", X"78", X"B1", X"20", X"FB", --7C80
  X"0B", X"78", X"B1", X"20", X"FB", X"18", X"D9", X"13", --7C88
  X"00", X"31", X"39", X"13", X"01", X"38", X"36", X"00", --7C90
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --7C98
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --7CA0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --7CA8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --7CB0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --7CB8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --7CC0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --7CC8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --7CD0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --7CD8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --7CE0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --7CE8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --7CF0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --7CF8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --7D00
  X"00", X"10", X"10", X"10", X"10", X"00", X"10", X"00", --7D08
  X"00", X"24", X"24", X"00", X"00", X"00", X"00", X"00", --7D10
  X"00", X"24", X"7E", X"24", X"24", X"7E", X"24", X"00", --7D18
  X"00", X"08", X"3E", X"28", X"3E", X"0A", X"3E", X"08", --7D20
  X"00", X"62", X"64", X"08", X"10", X"26", X"46", X"00", --7D28
  X"00", X"10", X"28", X"10", X"2A", X"44", X"3A", X"00", --7D30
  X"00", X"08", X"10", X"00", X"00", X"00", X"00", X"00", --7D38
  X"00", X"04", X"08", X"08", X"08", X"08", X"04", X"00", --7D40
  X"00", X"20", X"10", X"10", X"10", X"10", X"20", X"00", --7D48
  X"00", X"00", X"14", X"08", X"3E", X"08", X"14", X"00", --7D50
  X"00", X"00", X"08", X"08", X"3E", X"08", X"08", X"00", --7D58
  X"00", X"00", X"00", X"00", X"00", X"08", X"08", X"10", --7D60
  X"00", X"00", X"00", X"00", X"3E", X"00", X"00", X"00", --7D68
  X"00", X"00", X"00", X"00", X"00", X"18", X"18", X"00", --7D70
  X"00", X"00", X"02", X"04", X"08", X"10", X"20", X"00", --7D78
  X"00", X"3C", X"46", X"4A", X"52", X"62", X"3C", X"00", --7D80
  X"00", X"18", X"28", X"08", X"08", X"08", X"3E", X"00", --7D88
  X"00", X"3C", X"42", X"02", X"3C", X"40", X"7E", X"00", --7D90
  X"00", X"3C", X"42", X"0C", X"02", X"42", X"3C", X"00", --7D98
  X"00", X"08", X"18", X"28", X"48", X"7E", X"08", X"00", --7DA0
  X"00", X"7E", X"40", X"7C", X"02", X"42", X"3C", X"00", --7DA8
  X"00", X"3C", X"40", X"7C", X"42", X"42", X"3C", X"00", --7DB0
  X"00", X"7E", X"02", X"04", X"08", X"10", X"10", X"00", --7DB8
  X"00", X"3C", X"42", X"3C", X"42", X"42", X"3C", X"00", --7DC0
  X"00", X"3C", X"42", X"42", X"3E", X"02", X"3C", X"00", --7DC8
  X"00", X"00", X"00", X"10", X"00", X"00", X"10", X"00", --7DD0
  X"00", X"00", X"10", X"00", X"00", X"10", X"10", X"20", --7DD8
  X"00", X"00", X"04", X"08", X"10", X"08", X"04", X"00", --7DE0
  X"00", X"00", X"00", X"3E", X"00", X"3E", X"00", X"00", --7DE8
  X"00", X"00", X"10", X"08", X"04", X"08", X"10", X"00", --7DF0
  X"00", X"3C", X"42", X"04", X"08", X"00", X"08", X"00", --7DF8
  X"00", X"3C", X"4A", X"56", X"5E", X"40", X"3C", X"00", --7E00
  X"00", X"3C", X"42", X"42", X"7E", X"42", X"42", X"00", --7E08
  X"00", X"7C", X"42", X"7C", X"42", X"42", X"7C", X"00", --7E10
  X"00", X"3C", X"42", X"40", X"40", X"42", X"3C", X"00", --7E18
  X"00", X"78", X"44", X"42", X"42", X"44", X"78", X"00", --7E20
  X"00", X"7E", X"40", X"7C", X"40", X"40", X"7E", X"00", --7E28
  X"00", X"7E", X"40", X"7C", X"40", X"40", X"40", X"00", --7E30
  X"00", X"3C", X"42", X"40", X"4E", X"42", X"3C", X"00", --7E38
  X"00", X"42", X"42", X"7E", X"42", X"42", X"42", X"00", --7E40
  X"00", X"3E", X"08", X"08", X"08", X"08", X"3E", X"00", --7E48
  X"00", X"02", X"02", X"02", X"42", X"42", X"3C", X"00", --7E50
  X"00", X"44", X"48", X"70", X"48", X"44", X"42", X"00", --7E58
  X"00", X"40", X"40", X"40", X"40", X"40", X"7E", X"00", --7E60
  X"00", X"42", X"66", X"5A", X"42", X"42", X"42", X"00", --7E68
  X"00", X"42", X"62", X"52", X"4A", X"46", X"42", X"00", --7E70
  X"00", X"3C", X"42", X"42", X"42", X"42", X"3C", X"00", --7E78
  X"00", X"7C", X"42", X"42", X"7C", X"40", X"40", X"00", --7E80
  X"00", X"3C", X"42", X"42", X"52", X"4A", X"3C", X"00", --7E88
  X"00", X"7C", X"42", X"42", X"7C", X"44", X"42", X"00", --7E90
  X"00", X"3C", X"40", X"3C", X"02", X"42", X"3C", X"00", --7E98
  X"00", X"FE", X"10", X"10", X"10", X"10", X"10", X"00", --7EA0
  X"00", X"42", X"42", X"42", X"42", X"42", X"3C", X"00", --7EA8
  X"00", X"42", X"42", X"42", X"42", X"24", X"18", X"00", --7EB0
  X"00", X"42", X"42", X"42", X"42", X"5A", X"24", X"00", --7EB8
  X"00", X"42", X"24", X"18", X"18", X"24", X"42", X"00", --7EC0
  X"00", X"82", X"44", X"28", X"10", X"10", X"10", X"00", --7EC8
  X"00", X"7E", X"04", X"08", X"10", X"20", X"7E", X"00", --7ED0
  X"00", X"0E", X"08", X"08", X"08", X"08", X"0E", X"00", --7ED8
  X"00", X"00", X"40", X"20", X"10", X"08", X"04", X"00", --7EE0
  X"00", X"70", X"10", X"10", X"10", X"10", X"70", X"00", --7EE8
  X"00", X"10", X"38", X"54", X"10", X"10", X"10", X"00", --7EF0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"FF", --7EF8
  X"00", X"1C", X"22", X"78", X"20", X"20", X"7E", X"00", --7F00
  X"00", X"00", X"38", X"04", X"3C", X"44", X"3C", X"00", --7F08
  X"00", X"20", X"20", X"3C", X"22", X"22", X"3C", X"00", --7F10
  X"00", X"00", X"1C", X"20", X"20", X"20", X"1C", X"00", --7F18
  X"00", X"04", X"04", X"3C", X"44", X"44", X"3C", X"00", --7F20
  X"00", X"00", X"38", X"44", X"78", X"40", X"3C", X"00", --7F28
  X"00", X"0C", X"10", X"18", X"10", X"10", X"10", X"00", --7F30
  X"00", X"00", X"3C", X"44", X"44", X"3C", X"04", X"38", --7F38
  X"00", X"40", X"40", X"78", X"44", X"44", X"44", X"00", --7F40
  X"00", X"10", X"00", X"30", X"10", X"10", X"38", X"00", --7F48
  X"00", X"04", X"00", X"04", X"04", X"04", X"24", X"18", --7F50
  X"00", X"20", X"28", X"30", X"30", X"28", X"24", X"00", --7F58
  X"00", X"10", X"10", X"10", X"10", X"10", X"0C", X"00", --7F60
  X"00", X"00", X"68", X"54", X"54", X"54", X"54", X"00", --7F68
  X"00", X"00", X"78", X"44", X"44", X"44", X"44", X"00", --7F70
  X"00", X"00", X"38", X"44", X"44", X"44", X"38", X"00", --7F78
  X"00", X"00", X"78", X"44", X"44", X"78", X"40", X"40", --7F80
  X"00", X"00", X"3C", X"44", X"44", X"3C", X"04", X"06", --7F88
  X"00", X"00", X"1C", X"20", X"20", X"20", X"20", X"00", --7F90
  X"00", X"00", X"38", X"40", X"38", X"04", X"78", X"00", --7F98
  X"00", X"10", X"38", X"10", X"10", X"10", X"0C", X"00", --7FA0
  X"00", X"00", X"44", X"44", X"44", X"44", X"38", X"00", --7FA8
  X"00", X"00", X"44", X"44", X"28", X"28", X"10", X"00", --7FB0
  X"00", X"00", X"44", X"54", X"54", X"54", X"28", X"00", --7FB8
  X"00", X"00", X"44", X"28", X"10", X"28", X"44", X"00", --7FC0
  X"00", X"00", X"44", X"44", X"44", X"3C", X"04", X"38", --7FC8
  X"00", X"00", X"7C", X"08", X"10", X"20", X"7C", X"00", --7FD0
  X"00", X"0E", X"08", X"30", X"08", X"08", X"0E", X"00", --7FD8
  X"00", X"08", X"08", X"08", X"08", X"08", X"08", X"00", --7FE0
  X"00", X"70", X"10", X"0C", X"10", X"10", X"70", X"00", --7FE8
  X"00", X"14", X"28", X"00", X"00", X"00", X"00", X"00", --7FF0
  X"3C", X"42", X"99", X"A1", X"A1", X"99", X"42", X"3C");--7FF8

begin

  process (clk)
  begin
    if(rising_edge(clk)) then
      if wr='1' then
        ram(to_integer(unsigned(addr))) <= din;
      end if;
      dout <= ram(to_integer(unsigned(addr)));
    end if; 
  end process;

end architecture;
