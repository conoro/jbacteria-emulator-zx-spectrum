library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is port(
    clk   : in  std_logic;
    addr  : in  std_logic_vector(13 downto 0);
    dout  : out std_logic_vector(7 downto 0));
end rom;

architecture behavioral of rom is

  type rom_t is array (0 to 16383) of std_logic_vector(7 downto 0);
  signal rom : rom_t := (
  X"F3", X"3E", X"3F", X"ED", X"47", X"31", X"00", X"80", --0000
  X"00", X"00", X"00", X"00", X"00", X"00", X"21", X"3A", --0008
  X"01", X"22", X"1A", X"60", X"CD", X"1A", X"00", X"C3", --0010
  X"75", X"05", X"CD", X"18", X"02", X"06", X"1A", X"21", --0018
  X"00", X"60", X"36", X"00", X"23", X"10", X"FB", X"21", --0020
  X"D7", X"0A", X"22", X"00", X"60", X"3E", X"06", X"32", --0028
  X"02", X"60", X"CD", X"F0", X"00", X"21", X"B4", X"2D", --0030
  X"22", X"00", X"60", X"3E", X"1E", X"32", X"02", X"60", --0038
  X"CD", X"F0", X"00", X"3E", X"19", X"32", X"02", X"60", --0040
  X"CD", X"41", X"01", X"3E", X"1F", X"32", X"02", X"60", --0048
  X"CD", X"41", X"01", X"3E", X"26", X"32", X"02", X"60", --0050
  X"CD", X"41", X"01", X"3E", X"0C", X"32", X"9B", X"6E", --0058
  X"AF", X"32", X"9C", X"6E", X"3E", X"08", X"32", X"A1", --0060
  X"6E", X"3E", X"02", X"32", X"9F", X"6E", X"32", X"A0", --0068
  X"6E", X"21", X"C9", X"00", X"22", X"A2", X"6E", X"2A", --0070
  X"E6", X"00", X"22", X"9D", X"6E", X"CD", X"A1", X"17", --0078
  X"21", X"CF", X"00", X"22", X"A2", X"6E", X"2A", X"E8", --0080
  X"00", X"22", X"9D", X"6E", X"CD", X"A1", X"17", X"3E", --0088
  X"08", X"32", X"A1", X"6E", X"3E", X"04", X"32", X"9F", --0090
  X"6E", X"32", X"A0", X"6E", X"21", X"D8", X"00", X"22", --0098
  X"A2", X"6E", X"2A", X"EA", X"00", X"22", X"9D", X"6E", --00A0
  X"CD", X"A1", X"17", X"21", X"DE", X"00", X"22", X"A2", --00A8
  X"6E", X"2A", X"EC", X"00", X"22", X"9D", X"6E", X"CD", --00B0
  X"A1", X"17", X"06", X"0A", X"C5", X"01", X"FF", X"FF", --00B8
  X"0D", X"20", X"FD", X"10", X"FB", X"C1", X"10", X"F4", --00C0
  X"C9", X"50", X"53", X"49", X"4F", X"4E", X"FF", X"53", --00C8
  X"4F", X"46", X"54", X"57", X"41", X"52", X"45", X"FF", --00D0
  X"53", X"50", X"41", X"43", X"45", X"FF", X"52", X"41", --00D8
  X"49", X"44", X"45", X"52", X"53", X"FF", X"19", X"23", --00E0
  X"05", X"32", X"2A", X"64", X"16", X"87", X"C8", X"03", --00E8
  X"AF", X"CD", X"6A", X"13", X"21", X"00", X"03", X"22", --00F0
  X"04", X"60", X"2A", X"04", X"60", X"CD", X"67", X"17", --00F8
  X"ED", X"5B", X"02", X"60", X"CD", X"82", X"13", X"22", --0100
  X"06", X"60", X"2A", X"04", X"60", X"CD", X"9C", X"17", --0108
  X"ED", X"5B", X"02", X"60", X"CD", X"82", X"13", X"3A", --0110
  X"00", X"60", X"85", X"4F", X"3A", X"00", X"60", X"95", --0118
  X"6F", X"3A", X"06", X"60", X"47", X"3A", X"01", X"60", --0120
  X"80", X"47", X"60", X"CD", X"EC", X"12", X"ED", X"4B", --0128
  X"04", X"60", X"0B", X"0B", X"ED", X"43", X"04", X"60", --0130
  X"21", X"00", X"01", X"B7", X"ED", X"42", X"38", X"BA", --0138
  X"C9", X"21", X"00", X"04", X"22", X"04", X"60", X"3A", --0140
  X"02", X"60", X"CB", X"3F", X"32", X"0A", X"60", X"3A", --0148
  X"02", X"60", X"CB", X"27", X"32", X"08", X"60", X"2A", --0150
  X"EE", X"00", X"CD", X"67", X"17", X"32", X"0C", X"60", --0158
  X"ED", X"5B", X"08", X"60", X"CD", X"82", X"13", X"22", --0160
  X"0E", X"60", X"3A", X"0C", X"60", X"ED", X"5B", X"0A", --0168
  X"60", X"CD", X"82", X"13", X"22", X"10", X"60", X"2A", --0170
  X"EE", X"00", X"CD", X"9C", X"17", X"32", X"0D", X"60", --0178
  X"ED", X"5B", X"08", X"60", X"CD", X"82", X"13", X"22", --0180
  X"12", X"60", X"ED", X"5B", X"0A", X"60", X"3A", X"0D", --0188
  X"60", X"CD", X"82", X"13", X"22", X"14", X"60", X"2A", --0190
  X"04", X"60", X"CD", X"9C", X"17", X"ED", X"5B", X"12", --0198
  X"60", X"CD", X"82", X"13", X"22", X"16", X"60", X"2A", --01A0
  X"04", X"60", X"CD", X"67", X"17", X"ED", X"5B", X"10", --01A8
  X"60", X"CD", X"82", X"13", X"ED", X"4B", X"16", X"60", --01B0
  X"09", X"3A", X"00", X"60", X"85", X"32", X"16", X"60", --01B8
  X"2A", X"04", X"60", X"CD", X"67", X"17", X"ED", X"5B", --01C0
  X"14", X"60", X"CD", X"82", X"13", X"22", X"18", X"60", --01C8
  X"2A", X"04", X"60", X"CD", X"9C", X"17", X"ED", X"5B", --01D0
  X"0E", X"60", X"CD", X"82", X"13", X"ED", X"5B", X"18", --01D8
  X"60", X"EB", X"B7", X"ED", X"52", X"3A", X"01", X"60", --01E0
  X"85", X"47", X"3A", X"16", X"60", X"4F", X"ED", X"5B", --01E8
  X"04", X"60", X"B7", X"21", X"FE", X"01", X"ED", X"52", --01F0
  X"30", X"05", X"CD", X"42", X"14", X"18", X"03", X"CD", --01F8
  X"4F", X"14", X"ED", X"4B", X"04", X"60", X"0B", X"0B", --0200
  X"0B", X"0B", X"ED", X"43", X"04", X"60", X"21", X"00", --0208
  X"00", X"B7", X"ED", X"42", X"DA", X"97", X"01", X"C9", --0210
  X"CD", X"AD", X"12", X"3E", X"01", X"32", X"48", X"5C", --0218
  X"3E", X"01", X"D3", X"FE", X"3E", X"0E", X"57", X"5F", --0220
  X"21", X"00", X"00", X"39", X"31", X"00", X"5B", X"01", --0228
  X"80", X"01", X"D5", X"0B", X"79", X"B0", X"20", X"FA", --0230
  X"F9", X"C9", X"00", X"00", X"00", X"00", X"00", X"00", --0238
  X"00", X"00", X"00", X"10", X"10", X"10", X"10", X"00", --0240
  X"10", X"00", X"00", X"24", X"24", X"00", X"00", X"00", --0248
  X"00", X"00", X"00", X"24", X"7E", X"24", X"24", X"7E", --0250
  X"24", X"00", X"00", X"08", X"3E", X"28", X"3E", X"0A", --0258
  X"3E", X"08", X"00", X"62", X"64", X"08", X"10", X"26", --0260
  X"46", X"00", X"00", X"10", X"28", X"10", X"2A", X"44", --0268
  X"3A", X"00", X"00", X"08", X"10", X"00", X"00", X"00", --0270
  X"00", X"00", X"00", X"04", X"08", X"08", X"08", X"08", --0278
  X"04", X"00", X"00", X"20", X"10", X"10", X"10", X"10", --0280
  X"20", X"00", X"00", X"00", X"14", X"08", X"3E", X"08", --0288
  X"14", X"00", X"00", X"00", X"08", X"08", X"3E", X"08", --0290
  X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"08", --0298
  X"08", X"10", X"00", X"00", X"00", X"00", X"3E", X"00", --02A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"18", --02A8
  X"18", X"00", X"00", X"00", X"02", X"04", X"08", X"10", --02B0
  X"20", X"00", X"00", X"3C", X"46", X"4A", X"52", X"62", --02B8
  X"3C", X"00", X"00", X"18", X"28", X"08", X"08", X"08", --02C0
  X"3E", X"00", X"00", X"3C", X"42", X"02", X"3C", X"40", --02C8
  X"7E", X"00", X"00", X"3C", X"42", X"0C", X"02", X"42", --02D0
  X"3C", X"00", X"00", X"08", X"18", X"28", X"48", X"7E", --02D8
  X"08", X"00", X"00", X"7E", X"40", X"7C", X"02", X"42", --02E0
  X"3C", X"00", X"00", X"3C", X"40", X"7C", X"42", X"42", --02E8
  X"3C", X"00", X"00", X"7E", X"02", X"04", X"08", X"10", --02F0
  X"10", X"00", X"00", X"3C", X"42", X"3C", X"42", X"42", --02F8
  X"3C", X"00", X"00", X"3C", X"42", X"42", X"3E", X"02", --0300
  X"3C", X"00", X"00", X"00", X"00", X"10", X"00", X"00", --0308
  X"10", X"00", X"00", X"00", X"10", X"00", X"00", X"10", --0310
  X"10", X"20", X"00", X"00", X"04", X"08", X"10", X"08", --0318
  X"04", X"00", X"00", X"00", X"00", X"3E", X"00", X"3E", --0320
  X"00", X"00", X"00", X"00", X"10", X"08", X"04", X"08", --0328
  X"10", X"00", X"00", X"3C", X"42", X"04", X"08", X"00", --0330
  X"08", X"00", X"00", X"3C", X"4A", X"56", X"5E", X"40", --0338
  X"3C", X"00", X"00", X"3C", X"42", X"42", X"7E", X"42", --0340
  X"42", X"00", X"00", X"7C", X"42", X"7C", X"42", X"42", --0348
  X"7C", X"00", X"00", X"3C", X"42", X"40", X"40", X"42", --0350
  X"3C", X"00", X"00", X"78", X"44", X"42", X"42", X"44", --0358
  X"78", X"00", X"00", X"7E", X"40", X"7C", X"40", X"40", --0360
  X"7E", X"00", X"00", X"7E", X"40", X"7C", X"40", X"40", --0368
  X"40", X"00", X"00", X"3C", X"42", X"40", X"4E", X"42", --0370
  X"3C", X"00", X"00", X"42", X"42", X"7E", X"42", X"42", --0378
  X"42", X"00", X"00", X"3E", X"08", X"08", X"08", X"08", --0380
  X"3E", X"00", X"00", X"02", X"02", X"02", X"42", X"42", --0388
  X"3C", X"00", X"00", X"44", X"48", X"70", X"48", X"44", --0390
  X"42", X"00", X"00", X"40", X"40", X"40", X"40", X"40", --0398
  X"7E", X"00", X"00", X"42", X"66", X"5A", X"42", X"42", --03A0
  X"42", X"00", X"00", X"42", X"62", X"52", X"4A", X"46", --03A8
  X"42", X"00", X"00", X"3C", X"42", X"42", X"42", X"42", --03B0
  X"3C", X"00", X"00", X"7C", X"42", X"42", X"7C", X"40", --03B8
  X"40", X"00", X"00", X"3C", X"42", X"42", X"52", X"4A", --03C0
  X"3C", X"00", X"00", X"7C", X"42", X"42", X"7C", X"44", --03C8
  X"42", X"00", X"00", X"3C", X"40", X"3C", X"02", X"42", --03D0
  X"3C", X"00", X"00", X"FE", X"10", X"10", X"10", X"10", --03D8
  X"10", X"00", X"00", X"42", X"42", X"42", X"42", X"42", --03E0
  X"3C", X"00", X"00", X"42", X"42", X"42", X"42", X"24", --03E8
  X"18", X"00", X"00", X"42", X"42", X"42", X"42", X"5A", --03F0
  X"24", X"00", X"00", X"42", X"24", X"18", X"18", X"24", --03F8
  X"42", X"00", X"00", X"82", X"44", X"28", X"10", X"10", --0400
  X"10", X"00", X"00", X"7E", X"04", X"08", X"10", X"20", --0408
  X"7E", X"00", X"00", X"0E", X"08", X"08", X"08", X"08", --0410
  X"0E", X"00", X"00", X"00", X"40", X"20", X"10", X"08", --0418
  X"04", X"00", X"00", X"70", X"10", X"10", X"10", X"10", --0420
  X"70", X"00", X"00", X"10", X"38", X"54", X"10", X"10", --0428
  X"10", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0430
  X"00", X"FF", X"00", X"1C", X"22", X"78", X"20", X"20", --0438
  X"7E", X"00", X"00", X"00", X"38", X"04", X"3C", X"44", --0440
  X"3C", X"00", X"00", X"20", X"20", X"3C", X"22", X"22", --0448
  X"3C", X"00", X"00", X"00", X"1C", X"20", X"20", X"20", --0450
  X"1C", X"00", X"00", X"04", X"04", X"3C", X"44", X"44", --0458
  X"3C", X"00", X"00", X"00", X"38", X"44", X"78", X"40", --0460
  X"3C", X"00", X"00", X"0C", X"10", X"18", X"10", X"10", --0468
  X"10", X"00", X"00", X"00", X"3C", X"44", X"44", X"3C", --0470
  X"04", X"38", X"00", X"40", X"40", X"78", X"44", X"44", --0478
  X"44", X"00", X"00", X"10", X"00", X"30", X"10", X"10", --0480
  X"38", X"00", X"00", X"04", X"00", X"04", X"04", X"04", --0488
  X"24", X"18", X"00", X"20", X"28", X"30", X"30", X"28", --0490
  X"24", X"00", X"00", X"10", X"10", X"10", X"10", X"10", --0498
  X"0C", X"00", X"00", X"00", X"68", X"54", X"54", X"54", --04A0
  X"54", X"00", X"00", X"00", X"78", X"44", X"44", X"44", --04A8
  X"44", X"00", X"00", X"00", X"38", X"44", X"44", X"44", --04B0
  X"38", X"00", X"00", X"00", X"78", X"44", X"44", X"78", --04B8
  X"40", X"40", X"00", X"00", X"3C", X"44", X"44", X"3C", --04C0
  X"04", X"06", X"00", X"00", X"1C", X"20", X"20", X"20", --04C8
  X"20", X"00", X"00", X"00", X"38", X"40", X"38", X"04", --04D0
  X"78", X"00", X"00", X"10", X"38", X"10", X"10", X"10", --04D8
  X"0C", X"00", X"00", X"00", X"44", X"44", X"44", X"44", --04E0
  X"38", X"00", X"00", X"00", X"44", X"44", X"28", X"28", --04E8
  X"10", X"00", X"00", X"00", X"44", X"54", X"54", X"54", --04F0
  X"28", X"00", X"00", X"00", X"44", X"28", X"10", X"28", --04F8
  X"44", X"00", X"00", X"00", X"44", X"44", X"44", X"3C", --0500
  X"04", X"38", X"00", X"00", X"7C", X"08", X"10", X"20", --0508
  X"7C", X"00", X"00", X"0E", X"08", X"30", X"08", X"08", --0510
  X"0E", X"00", X"00", X"08", X"08", X"08", X"08", X"08", --0518
  X"08", X"00", X"00", X"70", X"10", X"0C", X"10", X"10", --0520
  X"70", X"00", X"00", X"14", X"28", X"00", X"00", X"00", --0528
  X"00", X"00", X"3C", X"42", X"99", X"A1", X"A1", X"99", --0530
  X"42", X"3C", X"05", X"06", X"04", X"04", X"02", X"02", --0538
  X"07", X"03", X"01", X"01", X"01", X"00", X"00", X"00", --0540
  X"03", X"05", X"00", X"00", X"37", X"0B", X"0B", X"0B", --0548
  X"0B", X"0B", X"05", X"05", X"05", X"05", X"05", X"05", --0550
  X"05", X"05", X"05", X"05", X"05", X"00", X"00", X"04", --0558
  X"01", X"00", X"0B", X"00", X"B8", X"00", X"00", X"00", --0560
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0568
  X"00", X"00", X"00", X"00", X"08", X"F3", X"31", X"00", --0570
  X"80", X"21", X"00", X"00", X"22", X"1E", X"60", X"22", --0578
  X"1C", X"60", X"21", X"35", X"82", X"22", X"A4", X"6E", --0580
  X"22", X"A6", X"6E", X"CD", X"01", X"06", X"CD", X"AD", --0588
  X"12", X"CD", X"AB", X"06", X"CD", X"D7", X"06", X"CD", --0590
  X"12", X"06", X"CD", X"F0", X"05", X"CD", X"8E", X"0E", --0598
  X"CD", X"99", X"07", X"CD", X"4E", X"0E", X"CD", X"E9", --05A0
  X"11", X"CD", X"8E", X"10", X"CD", X"1E", X"07", X"CD", --05A8
  X"13", X"07", X"CD", X"C1", X"0C", X"CD", X"BB", X"0A", --05B0
  X"3A", X"2A", X"60", X"B7", X"CA", X"66", X"06", X"CD", --05B8
  X"71", X"09", X"28", X"0A", X"3A", X"26", X"60", X"B7", --05C0
  X"CA", X"55", X"07", X"CD", X"D7", X"06", X"CD", X"6B", --05C8
  X"08", X"CD", X"E5", X"05", X"3A", X"26", X"60", X"B7", --05D0
  X"CA", X"55", X"07", X"3A", X"28", X"60", X"B7", X"C2", --05D8
  X"55", X"07", X"C3", X"33", X"06", X"3A", X"53", X"60", --05E0
  X"3D", X"32", X"53", X"60", X"C0", X"CD", X"B4", X"0F", --05E8
  X"3A", X"2A", X"60", X"CB", X"3F", X"CB", X"3F", X"47", --05F0
  X"CB", X"3F", X"80", X"C6", X"04", X"32", X"53", X"60", --05F8
  X"C9", X"3E", X"01", X"32", X"56", X"60", X"21", X"42", --0600
  X"05", X"11", X"20", X"60", X"01", X"0A", X"00", X"ED", --0608
  X"B0", X"C9", X"21", X"4C", X"05", X"11", X"2A", X"60", --0610
  X"01", X"29", X"00", X"ED", X"B0", X"3A", X"23", X"60", --0618
  X"3C", X"C8", X"32", X"23", X"60", X"FE", X"32", X"D0", --0620
  X"FE", X"09", X"D8", X"3A", X"27", X"60", X"3C", X"32", --0628
  X"27", X"60", X"C9", X"3A", X"50", X"60", X"B7", X"20", --0630
  X"06", X"3A", X"20", X"60", X"CD", X"5B", X"06", X"3A", --0638
  X"43", X"60", X"B7", X"20", X"06", X"3A", X"21", X"60", --0640
  X"CD", X"5B", X"06", X"3A", X"44", X"60", X"B7", X"C2", --0648
  X"AC", X"05", X"3A", X"22", X"60", X"CD", X"5B", X"06", --0650
  X"C3", X"AC", X"05", X"47", X"C5", X"06", X"00", X"00", --0658
  X"10", X"FD", X"C1", X"10", X"F7", X"C9", X"3A", X"29", --0660
  X"60", X"3C", X"FE", X"08", X"20", X"01", X"3D", X"32", --0668
  X"29", X"60", X"C3", X"97", X"05", X"32", X"54", X"60", --0670
  X"C5", X"CD", X"C6", X"12", X"3A", X"54", X"60", X"ED", --0678
  X"44", X"C6", X"05", X"28", X"05", X"DD", X"23", X"3D", --0680
  X"20", X"FB", X"DD", X"7E", X"00", X"DD", X"23", X"CD", --0688
  X"CB", X"13", X"C1", X"50", X"59", X"1C", X"D5", X"CD", --0690
  X"52", X"13", X"3A", X"54", X"60", X"3D", X"32", X"54", --0698
  X"60", X"20", X"E7", X"AF", X"CD", X"CB", X"13", X"C1", --06A0
  X"C3", X"52", X"13", X"ED", X"5B", X"1C", X"60", X"2A", --06A8
  X"1E", X"60", X"B7", X"ED", X"52", X"30", X"04", X"ED", --06B0
  X"53", X"1E", X"60", X"21", X"00", X"00", X"22", X"1C", --06B8
  X"60", X"CD", X"88", X"15", X"15", X"00", X"48", X"49", --06C0
  X"47", X"48", X"20", X"00", X"01", X"1A", X"00", X"2A", --06C8
  X"1E", X"60", X"3E", X"05", X"C3", X"75", X"06", X"11", --06D0
  X"00", X"40", X"CD", X"99", X"0A", X"3A", X"26", X"60", --06D8
  X"3D", X"28", X"2D", X"FA", X"10", X"07", X"32", X"55", --06E0
  X"60", X"ED", X"5B", X"41", X"60", X"D5", X"AF", X"32", --06E8
  X"42", X"60", X"3E", X"48", X"32", X"41", X"60", X"CD", --06F0
  X"4E", X"0E", X"3A", X"41", X"60", X"C6", X"18", X"32", --06F8
  X"41", X"60", X"3A", X"55", X"60", X"3D", X"32", X"55", --0700
  X"60", X"20", X"EC", X"D1", X"ED", X"53", X"41", X"60", --0708
  X"CD", X"C1", X"06", X"2A", X"1C", X"60", X"01", X"00", --0710
  X"00", X"3E", X"05", X"C3", X"75", X"06", X"3A", X"24", --0718
  X"60", X"B7", X"C0", X"2A", X"1C", X"60", X"01", X"64", --0720
  X"00", X"ED", X"42", X"D8", X"3E", X"01", X"32", X"24", --0728
  X"60", X"3A", X"26", X"60", X"3C", X"32", X"26", X"60", --0730
  X"06", X"08", X"3A", X"48", X"5C", X"C6", X"08", X"E6", --0738
  X"38", X"32", X"48", X"5C", X"CD", X"0D", X"16", X"0C", --0740
  X"28", X"12", X"1E", X"18", X"14", X"30", X"0A", X"00", --0748
  X"10", X"E8", X"C3", X"D7", X"06", X"CD", X"88", X"15", --0750
  X"00", X"17", X"47", X"41", X"4D", X"45", X"20", X"4F", --0758
  X"56", X"45", X"52", X"20", X"20", X"20", X"20", X"20", --0760
  X"20", X"20", X"48", X"49", X"54", X"20", X"46", X"49", --0768
  X"52", X"45", X"20", X"54", X"4F", X"20", X"50", X"4C", --0770
  X"41", X"59", X"00", X"06", X"19", X"CD", X"0D", X"16", --0778
  X"28", X"32", X"28", X"28", X"28", X"1E", X"28", X"14", --0780
  X"28", X"0A", X"00", X"10", X"F0", X"CD", X"D6", X"0C", --0788
  X"3A", X"4F", X"60", X"B7", X"28", X"F7", X"C3", X"8B", --0790
  X"05", X"3A", X"3A", X"05", X"E6", X"38", X"32", X"48", --0798
  X"5C", X"3A", X"3A", X"05", X"01", X"03", X"00", X"21", --07A0
  X"00", X"58", X"77", X"23", X"10", X"FC", X"0D", X"20", --07A8
  X"F9", X"CD", X"0D", X"16", X"64", X"64", X"00", X"01", --07B0
  X"00", X"01", X"3A", X"41", X"05", X"5F", X"16", X"20", --07B8
  X"CD", X"59", X"11", X"01", X"00", X"17", X"3A", X"40", --07C0
  X"05", X"5F", X"16", X"20", X"C3", X"59", X"11", X"13", --07C8
  X"01", X"14", X"02", X"03", X"03", X"07", X"03", X"0C", --07D0
  X"03", X"11", X"03", X"15", X"03", X"02", X"04", X"07", --07D8
  X"04", X"0C", X"04", X"11", X"04", X"16", X"04", X"03", --07E0
  X"05", X"07", X"05", X"0C", X"05", X"11", X"05", X"15", --07E8
  X"05", X"14", X"06", X"13", X"07", X"FF", X"03", X"01", --07F0
  X"02", X"02", X"01", X"03", X"05", X"03", X"0A", X"03", --07F8
  X"0F", X"03", X"13", X"03", X"00", X"04", X"05", X"04", --0800
  X"0A", X"04", X"0F", X"04", X"14", X"04", X"01", X"05", --0808
  X"05", X"05", X"0A", X"05", X"0F", X"05", X"13", X"05", --0810
  X"02", X"06", X"03", X"07", X"FF", X"04", X"01", X"03", --0818
  X"02", X"02", X"03", X"06", X"03", X"0B", X"03", X"10", --0820
  X"03", X"14", X"03", X"01", X"04", X"06", X"04", X"0B", --0828
  X"04", X"10", X"04", X"15", X"04", X"02", X"05", X"06", --0830
  X"05", X"0B", X"05", X"10", X"05", X"14", X"05", X"03", --0838
  X"06", X"04", X"07", X"FF", X"14", X"01", X"15", X"02", --0840
  X"04", X"03", X"08", X"03", X"0D", X"03", X"12", X"03", --0848
  X"16", X"03", X"03", X"04", X"08", X"04", X"0D", X"04", --0850
  X"12", X"04", X"17", X"04", X"04", X"05", X"08", X"05", --0858
  X"0D", X"05", X"12", X"05", X"16", X"05", X"15", X"06", --0860
  X"14", X"07", X"FF", X"3A", X"50", X"60", X"B7", X"20", --0868
  X"28", X"3A", X"A6", X"6E", X"FE", X"FF", X"C0", X"3A", --0870
  X"A7", X"6E", X"FE", X"19", X"D0", X"3A", X"A7", X"6E", --0878
  X"CB", X"47", X"28", X"0A", X"3E", X"01", X"32", X"50", --0880
  X"60", X"AF", X"32", X"51", X"60", X"C9", X"3E", X"FF", --0888
  X"32", X"50", X"60", X"3E", X"E9", X"32", X"51", X"60", --0890
  X"C9", X"3A", X"56", X"60", X"ED", X"44", X"32", X"56", --0898
  X"60", X"F2", X"25", X"09", X"DD", X"21", X"51", X"60", --08A0
  X"3A", X"50", X"60", X"FE", X"01", X"28", X"0E", X"21", --08A8
  X"CF", X"07", X"DD", X"35", X"00", X"AF", X"DD", X"BE", --08B0
  X"00", X"20", X"19", X"18", X"0D", X"21", X"1D", X"08", --08B8
  X"DD", X"34", X"00", X"3E", X"EA", X"DD", X"BE", X"00", --08C0
  X"20", X"0A", X"AF", X"32", X"50", X"60", X"11", X"20", --08C8
  X"40", X"C3", X"99", X"0A", X"3E", X"01", X"CD", X"2A", --08D0
  X"14", X"AF", X"CD", X"2A", X"14", X"3A", X"44", X"60", --08D8
  X"B7", X"C8", X"DD", X"21", X"45", X"60", X"DD", X"7E", --08E0
  X"01", X"FE", X"10", X"D0", X"3A", X"51", X"60", X"DD", --08E8
  X"BE", X"00", X"D0", X"C6", X"17", X"DD", X"BE", X"00", --08F0
  X"D8", X"CD", X"01", X"09", X"AF", X"32", X"50", X"60", --08F8
  X"C9", X"CD", X"CA", X"08", X"CD", X"34", X"09", X"CD", --0900
  X"0D", X"16", X"0A", X"FF", X"0A", X"C8", X"14", X"96", --0908
  X"05", X"C8", X"14", X"96", X"14", X"78", X"14", X"64", --0910
  X"14", X"50", X"14", X"3C", X"14", X"28", X"00", X"11", --0918
  X"20", X"40", X"C3", X"99", X"0A", X"CD", X"0D", X"16", --0920
  X"02", X"19", X"02", X"32", X"02", X"19", X"00", X"C9", --0928
  X"05", X"05", X"0A", X"14", X"3A", X"A7", X"6E", X"1F", --0930
  X"E6", X"03", X"21", X"30", X"09", X"CD", X"5F", X"09", --0938
  X"7E", X"47", X"2A", X"1C", X"60", X"CD", X"5F", X"09", --0940
  X"22", X"1C", X"60", X"3A", X"51", X"60", X"CB", X"3F", --0948
  X"CB", X"3F", X"CB", X"3F", X"4F", X"68", X"26", X"00", --0950
  X"06", X"01", X"3E", X"02", X"C3", X"75", X"06", X"85", --0958
  X"6F", X"D0", X"24", X"C9", X"00", X"00", X"00", X"01", --0960
  X"00", X"02", X"00", X"03", X"00", X"04", X"00", X"05", --0968
  X"FF", X"3E", X"04", X"32", X"5A", X"60", X"DD", X"21", --0970
  X"47", X"60", X"DD", X"7E", X"01", X"B7", X"28", X"05", --0978
  X"CD", X"02", X"0A", X"18", X"03", X"CD", X"9A", X"09", --0980
  X"CD", X"8E", X"09", X"20", X"ED", X"C9", X"DD", X"23", --0988
  X"DD", X"23", X"3A", X"5A", X"60", X"3D", X"32", X"5A", --0990
  X"60", X"C9", X"CD", X"B6", X"18", X"3A", X"A4", X"6E", --0998
  X"47", X"3A", X"27", X"60", X"B7", X"C8", X"B8", X"D8", --09A0
  X"3A", X"3D", X"60", X"32", X"57", X"60", X"3A", X"41", --09A8
  X"60", X"C6", X"07", X"47", X"3A", X"A6", X"6E", X"E6", --09B0
  X"0F", X"80", X"32", X"58", X"60", X"3A", X"A5", X"6E", --09B8
  X"FE", X"7F", X"30", X"06", X"3A", X"A6", X"6E", X"32", --09C0
  X"58", X"60", X"3A", X"57", X"60", X"DD", X"E5", X"CD", --09C8
  X"D1", X"0E", X"DD", X"7E", X"01", X"32", X"59", X"60", --09D0
  X"3A", X"58", X"60", X"CD", X"26", X"0B", X"DD", X"E1", --09D8
  X"20", X"0B", X"3A", X"57", X"60", X"3D", X"32", X"57", --09E0
  X"60", X"F2", X"CA", X"09", X"C9", X"3A", X"59", X"60", --09E8
  X"3C", X"3C", X"CB", X"27", X"CB", X"27", X"CB", X"27", --09F0
  X"DD", X"77", X"01", X"3A", X"58", X"60", X"DD", X"77", --09F8
  X"00", X"C9", X"21", X"64", X"09", X"3E", X"01", X"CD", --0A00
  X"2A", X"14", X"DD", X"7E", X"01", X"3C", X"FE", X"B9", --0A08
  X"D2", X"B6", X"0A", X"FE", X"B1", X"D2", X"32", X"0A", --0A10
  X"DD", X"77", X"01", X"C6", X"05", X"47", X"DD", X"4E", --0A18
  X"00", X"DD", X"E5", X"CD", X"42", X"12", X"DD", X"E1", --0A20
  X"C2", X"B6", X"0A", X"21", X"64", X"09", X"AF", X"C3", --0A28
  X"2A", X"14", X"DD", X"7E", X"00", X"47", X"3A", X"41", --0A30
  X"60", X"B8", X"30", X"53", X"C6", X"13", X"B8", X"38", --0A38
  X"4E", X"AF", X"32", X"41", X"60", X"06", X"08", X"3A", --0A40
  X"48", X"5C", X"C6", X"08", X"E6", X"38", X"32", X"48", --0A48
  X"5C", X"CD", X"0D", X"16", X"28", X"0A", X"28", X"14", --0A50
  X"28", X"28", X"28", X"50", X"00", X"10", X"E8", X"CD", --0A58
  X"96", X"0A", X"CD", X"0D", X"16", X"32", X"FF", X"FF", --0A60
  X"32", X"32", X"FF", X"00", X"3A", X"26", X"60", X"3D", --0A68
  X"32", X"26", X"60", X"C4", X"4E", X"0E", X"CD", X"7D", --0A70
  X"0A", X"F6", X"01", X"E1", X"C9", X"3E", X"04", X"32", --0A78
  X"5A", X"60", X"DD", X"21", X"47", X"60", X"CD", X"A9", --0A80
  X"0A", X"CD", X"8E", X"09", X"20", X"F8", X"C9", X"DD", --0A88
  X"7E", X"01", X"3C", X"C3", X"18", X"0A", X"11", X"E0", --0A90
  X"50", X"0E", X"08", X"AF", X"06", X"20", X"D5", X"12", --0A98
  X"13", X"10", X"FC", X"D1", X"14", X"0D", X"20", X"F4", --0AA0
  X"C9", X"DD", X"7E", X"01", X"B7", X"C8", X"21", X"64", --0AA8
  X"09", X"3E", X"01", X"CD", X"2A", X"14", X"DD", X"36", --0AB0
  X"01", X"00", X"C9", X"3A", X"44", X"60", X"B7", X"C8", --0AB8
  X"CD", X"C6", X"0A", X"C3", X"75", X"0C", X"3A", X"46", --0AC0
  X"60", X"CB", X"3F", X"CB", X"3F", X"CB", X"3F", X"3C", --0AC8
  X"32", X"5F", X"60", X"3A", X"3D", X"60", X"32", X"5D", --0AD0
  X"60", X"CD", X"D1", X"0E", X"3A", X"5F", X"60", X"DD", --0AD8
  X"BE", X"01", X"28", X"08", X"3A", X"5D", X"60", X"3D", --0AE0
  X"F2", X"D6", X"0A", X"C9", X"3A", X"45", X"60", X"CD", --0AE8
  X"26", X"0B", X"C8", X"C3", X"6D", X"0B", X"10", X"80", --0AF0
  X"09", X"10", X"49", X"20", X"26", X"40", X"10", X"80", --0AF8
  X"00", X"00", X"10", X"80", X"66", X"60", X"89", X"30", --0B00
  X"09", X"80", X"10", X"80", X"00", X"00", X"00", X"00", --0B08
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0B10
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0B18
  X"00", X"00", X"00", X"00", X"00", X"00", X"32", X"5B", --0B20
  X"60", X"CD", X"AE", X"10", X"DD", X"21", X"35", X"6E", --0B28
  X"3A", X"5B", X"60", X"47", X"CB", X"3F", X"CB", X"3F", --0B30
  X"CB", X"3F", X"32", X"5E", X"60", X"DD", X"96", X"04", --0B38
  X"38", X"29", X"CB", X"47", X"28", X"04", X"CB", X"50", --0B40
  X"20", X"21", X"DD", X"BE", X"05", X"30", X"1C", X"E6", --0B48
  X"FE", X"DD", X"86", X"04", X"32", X"5E", X"60", X"DD", --0B50
  X"96", X"02", X"32", X"5C", X"60", X"4F", X"06", X"00", --0B58
  X"DD", X"2A", X"35", X"6E", X"DD", X"09", X"DD", X"7E", --0B60
  X"02", X"B7", X"C9", X"AF", X"C9", X"CD", X"CC", X"0B", --0B68
  X"21", X"F6", X"0A", X"22", X"60", X"60", X"21", X"06", --0B70
  X"0B", X"22", X"62", X"60", X"CD", X"DD", X"0B", X"CD", --0B78
  X"3D", X"0E", X"CD", X"0D", X"16", X"10", X"50", X"20", --0B80
  X"28", X"40", X"14", X"80", X"0A", X"00", X"CD", X"5C", --0B88
  X"0C", X"21", X"16", X"0B", X"22", X"60", X"60", X"22", --0B90
  X"62", X"60", X"CD", X"DD", X"0B", X"3A", X"2A", X"60", --0B98
  X"3D", X"32", X"2A", X"60", X"C2", X"03", X"0C", X"CD", --0BA0
  X"7D", X"0A", X"06", X"28", X"3A", X"48", X"5C", X"C6", --0BA8
  X"08", X"E6", X"38", X"32", X"48", X"5C", X"CD", X"0D", --0BB0
  X"16", X"10", X"64", X"20", X"32", X"40", X"19", X"20", --0BB8
  X"32", X"00", X"10", X"E8", X"CD", X"CA", X"08", X"CD", --0BC0
  X"96", X"0A", X"E1", X"C9", X"06", X"20", X"11", X"16", --0BC8
  X"00", X"AF", X"DD", X"77", X"02", X"DD", X"77", X"03", --0BD0
  X"DD", X"19", X"10", X"F6", X"C9", X"ED", X"4B", X"5E", --0BD8
  X"60", X"CD", X"F8", X"15", X"2A", X"60", X"60", X"CD", --0BE0
  X"F5", X"0B", X"ED", X"4B", X"5E", X"60", X"04", X"CD", --0BE8
  X"F8", X"15", X"2A", X"62", X"60", X"06", X"08", X"ED", --0BF0
  X"A0", X"ED", X"A0", X"1B", X"1B", X"03", X"03", X"14", --0BF8
  X"10", X"F5", X"C9", X"21", X"2B", X"60", X"3A", X"5D", --0C00
  X"60", X"CD", X"70", X"0C", X"35", X"21", X"30", X"60", --0C08
  X"DD", X"21", X"35", X"6E", X"3A", X"5C", X"60", X"CB", --0C10
  X"3F", X"CD", X"70", X"0C", X"35", X"21", X"2B", X"60", --0C18
  X"3A", X"3D", X"60", X"3C", X"47", X"CD", X"70", X"0C", --0C20
  X"AF", X"2B", X"05", X"B6", X"28", X"FB", X"78", X"32", --0C28
  X"3D", X"60", X"06", X"FF", X"21", X"30", X"60", X"AF", --0C30
  X"2B", X"23", X"04", X"B6", X"28", X"FB", X"78", X"32", --0C38
  X"3F", X"60", X"21", X"30", X"60", X"3E", X"0B", X"47", --0C40
  X"04", X"CD", X"70", X"0C", X"AF", X"2B", X"05", X"B6", --0C48
  X"28", X"FB", X"78", X"32", X"40", X"60", X"C9", X"03", --0C50
  X"02", X"02", X"01", X"01", X"3A", X"5D", X"60", X"21", --0C58
  X"57", X"0C", X"CD", X"70", X"0C", X"7E", X"2A", X"1C", --0C60
  X"60", X"CD", X"70", X"0C", X"22", X"1C", X"60", X"C9", --0C68
  X"85", X"6F", X"D0", X"24", X"C9", X"DD", X"21", X"47", --0C70
  X"60", X"3E", X"04", X"32", X"64", X"60", X"ED", X"4B", --0C78
  X"45", X"60", X"DD", X"7E", X"01", X"B7", X"28", X"20", --0C80
  X"DD", X"7E", X"00", X"B9", X"20", X"1A", X"DD", X"7E", --0C88
  X"01", X"90", X"ED", X"44", X"FE", X"06", X"30", X"10", --0C90
  X"CD", X"A9", X"0A", X"CD", X"0D", X"16", X"04", X"18", --0C98
  X"08", X"0C", X"10", X"06", X"00", X"C3", X"3D", X"0E", --0CA0
  X"DD", X"23", X"DD", X"23", X"3A", X"64", X"60", X"3D", --0CA8
  X"32", X"64", X"60", X"20", X"CD", X"ED", X"4B", X"45", --0CB0
  X"60", X"05", X"CD", X"42", X"12", X"C8", X"C3", X"3D", --0CB8
  X"0E", X"CD", X"D6", X"0C", X"CD", X"2E", X"0D", X"3A", --0CC0
  X"44", X"60", X"B7", X"C2", X"1E", X"0E", X"3A", X"4F", --0CC8
  X"60", X"B7", X"C8", X"C3", X"FD", X"0D", X"01", X"FE", --0CD0
  X"FE", X"ED", X"58", X"01", X"FE", X"F7", X"ED", X"50", --0CD8
  X"3A", X"41", X"60", X"0E", X"00", X"CB", X"4B", X"28", --0CE0
  X"04", X"CB", X"42", X"20", X"04", X"B7", X"28", X"01", --0CE8
  X"0D", X"CB", X"53", X"28", X"04", X"CB", X"4A", X"20", --0CF0
  X"05", X"FE", X"EB", X"28", X"01", X"0C", X"79", X"32", --0CF8
  X"43", X"60", X"01", X"FE", X"7F", X"ED", X"58", X"CB", --0D00
  X"43", X"28", X"0E", X"CB", X"62", X"28", X"0A", X"3E", --0D08
  X"01", X"32", X"65", X"60", X"AF", X"32", X"4F", X"60", --0D10
  X"C9", X"CB", X"63", X"20", X"02", X"C1", X"C9", X"3A", --0D18
  X"65", X"60", X"B7", X"CA", X"14", X"0D", X"32", X"4F", --0D20
  X"60", X"AF", X"32", X"65", X"60", X"C9", X"3A", X"43", --0D28
  X"60", X"B7", X"C8", X"F2", X"37", X"0D", X"AF", X"DD", --0D30
  X"21", X"41", X"60", X"CD", X"53", X"0D", X"3E", X"01", --0D38
  X"CD", X"2A", X"14", X"AF", X"CD", X"2A", X"14", X"3A", --0D40
  X"43", X"60", X"47", X"3A", X"41", X"60", X"80", X"32", --0D48
  X"41", X"60", X"C9", X"21", X"5C", X"0D", X"B7", X"C0", --0D50
  X"21", X"A6", X"0D", X"C9", X"0A", X"00", X"09", X"01", --0D58
  X"01", X"02", X"09", X"02", X"13", X"02", X"01", X"03", --0D60
  X"09", X"03", X"13", X"03", X"01", X"04", X"06", X"04", --0D68
  X"12", X"04", X"01", X"05", X"01", X"06", X"06", X"06", --0D70
  X"12", X"06", X"01", X"07", X"07", X"07", X"13", X"07", --0D78
  X"FF", X"0B", X"00", X"0C", X"01", X"02", X"02", X"0C", --0D80
  X"02", X"14", X"02", X"02", X"03", X"0C", X"03", X"14", --0D88
  X"03", X"03", X"04", X"0F", X"04", X"14", X"04", X"14", --0D90
  X"05", X"03", X"06", X"0F", X"06", X"14", X"06", X"02", --0D98
  X"07", X"0E", X"07", X"14", X"07", X"FF", X"0A", X"00", --0DA0
  X"0B", X"01", X"01", X"02", X"0B", X"02", X"13", X"02", --0DA8
  X"01", X"03", X"0B", X"03", X"13", X"03", X"02", X"04", --0DB0
  X"0E", X"04", X"13", X"04", X"13", X"05", X"02", X"06", --0DB8
  X"0E", X"06", X"13", X"06", X"01", X"07", X"0D", X"07", --0DC0
  X"13", X"07", X"FF", X"09", X"00", X"08", X"01", X"00", --0DC8
  X"02", X"08", X"02", X"12", X"02", X"00", X"03", X"08", --0DD0
  X"03", X"12", X"03", X"00", X"04", X"05", X"04", X"11", --0DD8
  X"04", X"00", X"05", X"00", X"06", X"05", X"06", X"11", --0DE0
  X"06", X"00", X"07", X"06", X"07", X"12", X"07", X"FF", --0DE8
  X"00", X"00", X"00", X"01", X"00", X"02", X"00", X"03", --0DF0
  X"00", X"04", X"00", X"05", X"FF", X"CD", X"0D", X"16", --0DF8
  X"14", X"32", X"0A", X"64", X"05", X"C8", X"00", X"3E", --0E00
  X"01", X"32", X"44", X"60", X"3A", X"41", X"60", X"DD", --0E08
  X"21", X"45", X"60", X"C6", X"0A", X"DD", X"77", X"00", --0E10
  X"DD", X"36", X"01", X"B0", X"18", X"18", X"DD", X"21", --0E18
  X"45", X"60", X"21", X"F0", X"0D", X"3E", X"01", X"CD", --0E20
  X"2A", X"14", X"DD", X"7E", X"01", X"D6", X"04", X"FE", --0E28
  X"04", X"28", X"16", X"DD", X"77", X"01", X"21", X"F0", --0E30
  X"0D", X"AF", X"C3", X"2A", X"14", X"DD", X"21", X"45", --0E38
  X"60", X"21", X"F0", X"0D", X"3E", X"01", X"CD", X"2A", --0E40
  X"14", X"AF", X"32", X"44", X"60", X"C9", X"DD", X"E5", --0E48
  X"E5", X"3E", X"FF", X"32", X"43", X"60", X"3A", X"41", --0E50
  X"60", X"32", X"66", X"60", X"C6", X"28", X"32", X"41", --0E58
  X"60", X"CD", X"2E", X"0D", X"CD", X"0D", X"16", X"01", --0E60
  X"0F", X"00", X"3A", X"66", X"60", X"DD", X"BE", X"00", --0E68
  X"20", X"EF", X"E1", X"DD", X"E1", X"C9", X"0E", X"20", --0E70
  X"5E", X"23", X"56", X"23", X"06", X"0B", X"DD", X"73", --0E78
  X"00", X"DD", X"23", X"DD", X"72", X"00", X"DD", X"23", --0E80
  X"10", X"F4", X"0D", X"20", X"EB", X"C9", X"3A", X"29", --0E88
  X"60", X"C6", X"03", X"32", X"6A", X"60", X"21", X"AF", --0E90
  X"0F", X"22", X"68", X"60", X"3E", X"04", X"32", X"67", --0E98
  X"60", X"DD", X"21", X"6B", X"60", X"DD", X"36", X"00", --0EA0
  X"05", X"DD", X"23", X"3A", X"6A", X"60", X"DD", X"77", --0EA8
  X"00", X"DD", X"23", X"3C", X"3C", X"32", X"6A", X"60", --0EB0
  X"2A", X"68", X"60", X"7E", X"23", X"22", X"68", X"60", --0EB8
  X"CD", X"E2", X"0E", X"CD", X"76", X"0E", X"3A", X"67", --0EC0
  X"60", X"3D", X"32", X"67", X"60", X"F2", X"A5", X"0E", --0EC8
  X"C9", X"DD", X"21", X"6B", X"60", X"B7", X"C8", X"C5", --0ED0
  X"01", X"C2", X"02", X"DD", X"09", X"3D", X"20", X"FB", --0ED8
  X"C1", X"C9", X"21", X"EF", X"0E", X"B7", X"C8", X"01", --0EE0
  X"40", X"00", X"09", X"3D", X"20", X"FC", X"C9", X"1F", --0EE8
  X"80", X"3F", X"C0", X"7F", X"E0", X"FF", X"F0", X"DE", --0EF0
  X"F0", X"DE", X"F0", X"DE", X"F0", X"FF", X"F0", X"3F", --0EF8
  X"80", X"30", X"C0", X"60", X"60", X"C0", X"30", X"00", --0F00
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"1F", --0F08
  X"80", X"3F", X"C0", X"7F", X"E0", X"FF", X"F0", X"F7", --0F10
  X"B0", X"F7", X"B0", X"F7", X"B0", X"FF", X"F0", X"1F", --0F18
  X"80", X"19", X"80", X"19", X"80", X"19", X"80", X"00", --0F20
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C0", --0F28
  X"30", X"C0", X"30", X"FF", X"F0", X"86", X"10", X"E7", --0F30
  X"90", X"86", X"10", X"FF", X"F0", X"2F", X"40", X"4F", --0F38
  X"20", X"86", X"10", X"40", X"20", X"20", X"40", X"00", --0F40
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C0", --0F48
  X"30", X"C0", X"30", X"FF", X"F0", X"86", X"10", X"9E", --0F50
  X"70", X"86", X"10", X"FF", X"F0", X"2F", X"40", X"2F", --0F58
  X"40", X"26", X"40", X"20", X"40", X"20", X"40", X"00", --0F60
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"30", --0F68
  X"C0", X"30", X"C0", X"09", X"00", X"0F", X"00", X"1F", --0F70
  X"80", X"3F", X"C0", X"7F", X"E0", X"B0", X"D0", X"9F", --0F78
  X"90", X"09", X"00", X"10", X"80", X"09", X"00", X"00", --0F80
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C0", --0F88
  X"30", X"C0", X"30", X"20", X"40", X"16", X"80", X"1F", --0F90
  X"80", X"3F", X"C0", X"FF", X"F0", X"30", X"C0", X"1F", --0F98
  X"80", X"09", X"00", X"10", X"80", X"20", X"40", X"00", --0FA0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"02", --0FA8
  X"01", X"01", X"00", X"00", X"3A", X"3B", X"60", X"47", --0FB0
  X"3A", X"3D", X"60", X"B8", X"30", X"15", X"32", X"3B", --0FB8
  X"60", X"3A", X"3C", X"60", X"B7", X"20", X"0C", X"3A", --0FC0
  X"3B", X"60", X"CD", X"D1", X"0E", X"CD", X"AE", X"10", --0FC8
  X"CD", X"1A", X"10", X"3A", X"3B", X"60", X"B7", X"20", --0FD0
  X"06", X"CD", X"0D", X"16", X"0A", X"FA", X"00", X"CD", --0FD8
  X"D1", X"0E", X"CD", X"AE", X"10", X"3A", X"3C", X"60", --0FE0
  X"B7", X"28", X"1A", X"CD", X"3E", X"10", X"3A", X"3B", --0FE8
  X"60", X"B7", X"20", X"0C", X"32", X"3C", X"60", X"3A", --0FF0
  X"3E", X"60", X"ED", X"44", X"32", X"3E", X"60", X"C9", --0FF8
  X"3D", X"32", X"3B", X"60", X"C9", X"CD", X"83", X"10", --1000
  X"3A", X"3B", X"60", X"47", X"3A", X"3D", X"60", X"B8", --1008
  X"28", X"08", X"3A", X"3B", X"60", X"3C", X"32", X"3B", --1010
  X"60", X"C9", X"3A", X"3E", X"60", X"FE", X"01", X"28", --1018
  X"0C", X"3A", X"39", X"6E", X"B7", X"20", X"12", X"3E", --1020
  X"01", X"32", X"3C", X"60", X"C9", X"3A", X"39", X"6E", --1028
  X"47", X"3A", X"3A", X"6E", X"80", X"FE", X"20", X"28", --1030
  X"EE", X"AF", X"32", X"3B", X"60", X"C9", X"CD", X"0D", --1038
  X"16", X"08", X"FA", X"00", X"3A", X"38", X"6E", X"FE", --1040
  X"12", X"D4", X"7E", X"11", X"3A", X"38", X"6E", X"FE", --1048
  X"15", X"28", X"1E", X"47", X"0E", X"00", X"CD", X"F8", --1050
  X"15", X"CD", X"99", X"0A", X"ED", X"4B", X"37", X"6E", --1058
  X"04", X"DD", X"2A", X"35", X"6E", X"DD", X"71", X"00", --1060
  X"DD", X"70", X"01", X"CD", X"AE", X"10", X"C3", X"FD", --1068
  X"10", X"3E", X"01", X"32", X"28", X"60", X"CD", X"0D", --1070
  X"16", X"FA", X"64", X"FA", X"C8", X"FA", X"FA", X"FA", --1078
  X"FA", X"00", X"C9", X"ED", X"4B", X"37", X"6E", X"3A", --1080
  X"3E", X"60", X"81", X"4F", X"18", X"D3", X"3E", X"04", --1088
  X"32", X"3B", X"60", X"CD", X"D1", X"0E", X"CD", X"AE", --1090
  X"10", X"CD", X"FD", X"10", X"CD", X"0D", X"16", X"19", --1098
  X"F0", X"64", X"78", X"19", X"F0", X"00", X"3A", X"3B", --10A0
  X"60", X"3D", X"F2", X"90", X"10", X"C9", X"DD", X"22", --10A8
  X"35", X"6E", X"DD", X"4E", X"00", X"DD", X"46", X"01", --10B0
  X"ED", X"43", X"37", X"6E", X"3A", X"3F", X"60", X"3C", --10B8
  X"CB", X"27", X"4F", X"06", X"00", X"DD", X"09", X"3A", --10C0
  X"37", X"6E", X"1F", X"30", X"05", X"01", X"60", X"01", --10C8
  X"DD", X"09", X"DD", X"22", X"3C", X"6E", X"3A", X"37", --10D0
  X"6E", X"47", X"3A", X"3F", X"60", X"CB", X"27", X"80", --10D8
  X"32", X"39", X"6E", X"3A", X"3F", X"60", X"47", X"3A", --10E0
  X"40", X"60", X"90", X"CB", X"27", X"32", X"3A", X"6E", --10E8
  X"47", X"3A", X"39", X"6E", X"80", X"D6", X"20", X"ED", --10F0
  X"44", X"32", X"3B", X"6E", X"C9", X"CD", X"66", X"11", --10F8
  X"ED", X"4B", X"37", X"6E", X"CD", X"0C", X"11", X"ED", --1100
  X"4B", X"37", X"6E", X"04", X"3E", X"08", X"32", X"40", --1108
  X"6E", X"0E", X"00", X"CD", X"F8", X"15", X"ED", X"53", --1110
  X"3E", X"6E", X"CD", X"38", X"11", X"2A", X"3C", X"6E", --1118
  X"01", X"16", X"00", X"09", X"22", X"3C", X"6E", X"2A", --1120
  X"3E", X"6E", X"24", X"22", X"3E", X"6E", X"3A", X"40", --1128
  X"6E", X"3D", X"32", X"40", X"6E", X"20", X"E3", X"C9", --1130
  X"ED", X"5B", X"3E", X"6E", X"3A", X"39", X"6E", X"CD", --1138
  X"50", X"11", X"2A", X"3C", X"6E", X"ED", X"4B", X"3A", --1140
  X"6E", X"06", X"00", X"ED", X"B0", X"3A", X"3B", X"6E", --1148
  X"B7", X"C8", X"47", X"AF", X"12", X"13", X"10", X"FC", --1150
  X"C9", X"CD", X"41", X"13", X"3E", X"F8", X"A6", X"B3", --1158
  X"77", X"23", X"15", X"20", X"F7", X"C9", X"ED", X"4B", --1160
  X"37", X"6E", X"0E", X"00", X"21", X"3B", X"05", X"3A", --1168
  X"3B", X"60", X"85", X"6F", X"30", X"01", X"24", X"7E", --1170
  X"5F", X"16", X"40", X"C3", X"59", X"11", X"3A", X"25", --1178
  X"60", X"B7", X"C8", X"11", X"80", X"50", X"CD", X"99", --1180
  X"0A", X"11", X"A0", X"50", X"CD", X"99", X"0A", X"11", --1188
  X"C0", X"50", X"CD", X"99", X"0A", X"AF", X"32", X"25", --1190
  X"60", X"CD", X"0D", X"16", X"C8", X"0A", X"0A", X"C8", --1198
  X"C8", X"0A", X"0A", X"C8", X"C8", X"0A", X"32", X"FA", --11A0
  X"00", X"C9", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --11A8
  X"FF", X"FF", X"03", X"0F", X"1F", X"3F", X"7F", X"7F", --11B0
  X"FF", X"FF", X"C0", X"F0", X"F8", X"FC", X"FE", X"FE", --11B8
  X"FF", X"FF", X"FC", X"F0", X"E0", X"C0", X"80", X"80", --11C0
  X"00", X"00", X"3F", X"0F", X"07", X"03", X"01", X"01", --11C8
  X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --11D0
  X"00", X"00", X"31", X"30", X"30", X"32", X"00", X"30", --11D8
  X"30", X"30", X"30", X"00", X"35", X"33", X"34", X"35", --11E0
  X"00", X"3A", X"25", X"60", X"B7", X"C0", X"2A", X"1A", --11E8
  X"60", X"E5", X"21", X"2A", X"10", X"22", X"1A", X"60", --11F0
  X"3E", X"03", X"32", X"41", X"6E", X"01", X"05", X"14", --11F8
  X"21", X"DA", X"11", X"C5", X"3E", X"03", X"32", X"42", --1200
  X"6E", X"CD", X"91", X"15", X"0D", X"0D", X"0D", X"0D", --1208
  X"04", X"3A", X"42", X"6E", X"3D", X"32", X"42", X"6E", --1210
  X"20", X"EF", X"C1", X"79", X"C6", X"09", X"4F", X"3A", --1218
  X"41", X"6E", X"3D", X"32", X"41", X"6E", X"20", X"D8", --1220
  X"E1", X"22", X"1A", X"60", X"3E", X"01", X"32", X"25", --1228
  X"60", X"C9", X"FE", X"00", X"FF", X"00", X"01", X"00", --1230
  X"02", X"00", X"FF", X"FF", X"01", X"FF", X"FF", X"01", --1238
  X"01", X"01", X"3A", X"25", X"60", X"B7", X"C8", X"ED", --1240
  X"43", X"43", X"6E", X"78", X"FE", X"A2", X"38", X"5B", --1248
  X"FE", X"B8", X"30", X"57", X"CD", X"55", X"14", X"C8", --1250
  X"CD", X"B6", X"18", X"DD", X"21", X"32", X"12", X"3E", --1258
  X"08", X"32", X"41", X"6E", X"3A", X"43", X"6E", X"DD", --1260
  X"86", X"00", X"4F", X"3A", X"44", X"6E", X"DD", X"86", --1268
  X"01", X"47", X"DD", X"23", X"DD", X"23", X"3A", X"A4", --1270
  X"6E", X"17", X"32", X"A4", X"6E", X"DC", X"48", X"14", --1278
  X"3A", X"41", X"6E", X"3D", X"32", X"41", X"6E", X"20", --1280
  X"DB", X"ED", X"4B", X"43", X"6E", X"CD", X"48", X"14", --1288
  X"ED", X"4B", X"43", X"6E", X"04", X"CD", X"48", X"14", --1290
  X"ED", X"4B", X"43", X"6E", X"05", X"CD", X"48", X"14", --1298
  X"CD", X"0D", X"16", X"04", X"14", X"04", X"1E", X"00", --12A0
  X"F6", X"01", X"C9", X"AF", X"C9", X"21", X"00", X"40", --12A8
  X"0E", X"18", X"AF", X"47", X"77", X"23", X"10", X"FC", --12B0
  X"0D", X"20", X"F9", X"C9", X"10", X"27", X"E8", X"03", --12B8
  X"64", X"00", X"0A", X"00", X"01", X"00", X"DD", X"21", --12C0
  X"45", X"6E", X"06", X"05", X"ED", X"73", X"4A", X"6E", --12C8
  X"31", X"BC", X"12", X"D1", X"F6", X"FF", X"ED", X"52", --12D0
  X"3C", X"30", X"FB", X"19", X"DD", X"77", X"00", X"DD", --12D8
  X"23", X"10", X"F0", X"DD", X"21", X"45", X"6E", X"ED", --12E0
  X"7B", X"4A", X"6E", X"C9", X"11", X"01", X"01", X"22", --12E8
  X"4C", X"6E", X"79", X"95", X"D2", X"FB", X"12", X"1E", --12F0
  X"FF", X"ED", X"44", X"4F", X"78", X"94", X"D2", X"05", --12F8
  X"13", X"16", X"FF", X"ED", X"44", X"47", X"79", X"B8", --1300
  X"30", X"06", X"69", X"D5", X"AF", X"5F", X"18", X"07", --1308
  X"B1", X"C8", X"68", X"41", X"D5", X"16", X"00", X"60", --1310
  X"78", X"1F", X"85", X"38", X"03", X"BC", X"38", X"07", --1318
  X"94", X"4F", X"D9", X"C1", X"C5", X"18", X"04", X"4F", --1320
  X"D5", X"D9", X"C1", X"2A", X"4C", X"6E", X"78", X"84", --1328
  X"47", X"79", X"85", X"4F", X"ED", X"43", X"4C", X"6E", --1330
  X"CD", X"5E", X"13", X"D9", X"79", X"10", X"DB", X"D1", --1338
  X"C9", X"78", X"F6", X"C0", X"6F", X"26", X"02", X"29", --1340
  X"29", X"29", X"29", X"29", X"79", X"85", X"6F", X"D0", --1348
  X"24", X"C9", X"CD", X"F8", X"15", X"06", X"08", X"7E", --1350
  X"23", X"12", X"14", X"10", X"FA", X"C9", X"2A", X"4E", --1358
  X"6E", X"E9", X"42", X"14", X"48", X"14", X"4F", X"14", --1360
  X"55", X"14", X"E5", X"C5", X"E6", X"03", X"6F", X"26", --1368
  X"00", X"29", X"01", X"62", X"13", X"09", X"01", X"4E", --1370
  X"6E", X"7E", X"02", X"23", X"03", X"7E", X"02", X"C1", --1378
  X"E1", X"C9", X"A7", X"F2", X"8F", X"13", X"21", X"00", --1380
  X"00", X"B7", X"ED", X"52", X"EB", X"ED", X"44", X"4B", --1388
  X"5A", X"16", X"00", X"47", X"CB", X"7B", X"28", X"01", --1390
  X"15", X"62", X"CB", X"21", X"CB", X"13", X"CB", X"12", --1398
  X"79", X"CB", X"17", X"7B", X"6A", X"CB", X"17", X"CB", --13A0
  X"15", X"CB", X"14", X"81", X"4F", X"ED", X"5A", X"EB", --13A8
  X"21", X"00", X"00", X"78", X"06", X"07", X"CB", X"1F", --13B0
  X"30", X"08", X"19", X"CB", X"21", X"30", X"05", X"23", --13B8
  X"18", X"02", X"CB", X"21", X"CB", X"13", X"CB", X"12", --13C0
  X"10", X"EC", X"C9", X"21", X"DA", X"13", X"CB", X"27", --13C8
  X"CB", X"27", X"CB", X"27", X"85", X"6F", X"30", X"01", --13D0
  X"24", X"C9", X"7E", X"7E", X"66", X"66", X"66", X"66", --13D8
  X"7E", X"7E", X"18", X"18", X"18", X"18", X"18", X"18", --13E0
  X"18", X"18", X"7E", X"7E", X"06", X"7E", X"7E", X"60", --13E8
  X"7E", X"7E", X"7E", X"7E", X"06", X"7E", X"7E", X"06", --13F0
  X"7E", X"7E", X"60", X"60", X"6C", X"6C", X"7E", X"7E", --13F8
  X"0C", X"0C", X"7E", X"7E", X"60", X"7E", X"7E", X"06", --1400
  X"7E", X"7E", X"7E", X"7E", X"60", X"7E", X"7E", X"66", --1408
  X"7E", X"7E", X"7E", X"7E", X"06", X"06", X"06", X"06", --1410
  X"06", X"06", X"7E", X"7E", X"66", X"7E", X"7E", X"66", --1418
  X"7E", X"7E", X"7E", X"7E", X"66", X"7E", X"7E", X"06", --1420
  X"7E", X"7E", X"CD", X"6A", X"13", X"7E", X"23", X"B7", --1428
  X"F8", X"DD", X"86", X"00", X"4F", X"7E", X"23", X"DD", --1430
  X"86", X"01", X"47", X"E5", X"CD", X"5E", X"13", X"E1", --1438
  X"18", X"EB", X"CD", X"62", X"15", X"B6", X"77", X"C9", --1440
  X"CD", X"62", X"15", X"2F", X"A6", X"77", X"C9", X"CD", --1448
  X"62", X"15", X"AE", X"77", X"C9", X"CD", X"62", X"15", --1450
  X"A6", X"C9", X"80", X"40", X"20", X"10", X"08", X"04", --1458
  X"02", X"01", X"00", X"08", X"10", X"18", X"20", X"28", --1460
  X"30", X"38", X"01", X"09", X"11", X"19", X"21", X"29", --1468
  X"31", X"39", X"02", X"0A", X"12", X"1A", X"22", X"2A", --1470
  X"32", X"3A", X"03", X"0B", X"13", X"1B", X"23", X"2B", --1478
  X"33", X"3B", X"04", X"0C", X"14", X"1C", X"24", X"2C", --1480
  X"34", X"3C", X"05", X"0D", X"15", X"1D", X"25", X"2D", --1488
  X"35", X"3D", X"06", X"0E", X"16", X"1E", X"26", X"2E", --1490
  X"36", X"3E", X"07", X"0F", X"17", X"1F", X"27", X"2F", --1498
  X"37", X"3F", X"40", X"48", X"50", X"58", X"60", X"68", --14A0
  X"70", X"78", X"41", X"49", X"51", X"59", X"61", X"69", --14A8
  X"71", X"79", X"42", X"4A", X"52", X"5A", X"62", X"6A", --14B0
  X"72", X"7A", X"43", X"4B", X"53", X"5B", X"63", X"6B", --14B8
  X"73", X"7B", X"44", X"4C", X"54", X"5C", X"64", X"6C", --14C0
  X"74", X"7C", X"45", X"4D", X"55", X"5D", X"65", X"6D", --14C8
  X"75", X"7D", X"46", X"4E", X"56", X"5E", X"66", X"6E", --14D0
  X"76", X"7E", X"47", X"4F", X"57", X"5F", X"67", X"6F", --14D8
  X"77", X"7F", X"80", X"88", X"90", X"98", X"A0", X"A8", --14E0
  X"B0", X"B8", X"81", X"89", X"91", X"99", X"A1", X"A9", --14E8
  X"B1", X"B9", X"82", X"8A", X"92", X"9A", X"A2", X"AA", --14F0
  X"B2", X"BA", X"83", X"8B", X"93", X"9B", X"A3", X"AB", --14F8
  X"B3", X"BB", X"84", X"8C", X"94", X"9C", X"A4", X"AC", --1500
  X"B4", X"BC", X"85", X"8D", X"95", X"9D", X"A5", X"AD", --1508
  X"B5", X"BD", X"86", X"8E", X"96", X"9E", X"A6", X"AE", --1510
  X"B6", X"BE", X"87", X"8F", X"97", X"9F", X"A7", X"AF", --1518
  X"B7", X"BF", X"00", X"08", X"10", X"18", X"20", X"28", --1520
  X"30", X"38", X"01", X"09", X"11", X"19", X"21", X"29", --1528
  X"31", X"39", X"02", X"0A", X"12", X"1A", X"22", X"2A", --1530
  X"32", X"3A", X"03", X"0B", X"13", X"1B", X"23", X"2B", --1538
  X"33", X"3B", X"84", X"8C", X"94", X"9C", X"A4", X"AC", --1540
  X"B4", X"BC", X"85", X"8D", X"95", X"9D", X"A5", X"AD", --1548
  X"B5", X"BD", X"86", X"8E", X"96", X"9E", X"A6", X"AE", --1550
  X"B6", X"BE", X"87", X"8F", X"97", X"9F", X"A7", X"AF", --1558
  X"B7", X"BF", X"21", X"62", X"14", X"58", X"16", X"00", --1560
  X"19", X"66", X"69", X"A7", X"CB", X"1C", X"CB", X"1D", --1568
  X"37", X"CB", X"1C", X"CB", X"1D", X"A7", X"CB", X"1C", --1570
  X"CB", X"1D", X"EB", X"21", X"5A", X"14", X"79", X"E6", --1578
  X"07", X"4F", X"06", X"00", X"09", X"7E", X"EB", X"C9", --1580
  X"E1", X"CD", X"8D", X"15", X"E9", X"4E", X"23", X"46", --1588
  X"23", X"7E", X"23", X"B7", X"C8", X"FE", X"01", X"28", --1590
  X"F4", X"C5", X"E5", X"CD", X"EB", X"18", X"CD", X"52", --1598
  X"13", X"E1", X"C1", X"CD", X"A8", X"15", X"18", X"E9", --15A0
  X"0C", X"79", X"FE", X"20", X"C0", X"0E", X"00", X"04", --15A8
  X"78", X"FE", X"18", X"C0", X"06", X"00", X"C9", X"E1", --15B0
  X"ED", X"73", X"50", X"6E", X"31", X"85", X"6E", X"E5", --15B8
  X"FD", X"22", X"86", X"6E", X"D9", X"22", X"88", X"6E", --15C0
  X"ED", X"53", X"8A", X"6E", X"ED", X"43", X"8C", X"6E", --15C8
  X"D9", X"C9", X"ED", X"73", X"52", X"6E", X"ED", X"7B", --15D0
  X"50", X"6E", X"D9", X"2A", X"88", X"6E", X"ED", X"5B", --15D8
  X"8A", X"6E", X"ED", X"4B", X"8C", X"6E", X"D9", X"FD", --15E0
  X"2A", X"86", X"6E", X"FB", X"C9", X"ED", X"73", X"50", --15E8
  X"6E", X"ED", X"7B", X"52", X"6E", X"C3", X"C4", X"15", --15F0
  X"50", X"AF", X"CB", X"18", X"1F", X"CB", X"18", X"1F", --15F8
  X"CB", X"18", X"1F", X"B1", X"5F", X"42", X"3E", X"18", --1600
  X"A2", X"F6", X"40", X"57", X"C9", X"ED", X"53", X"8E", --1608
  X"6E", X"D1", X"C5", X"F5", X"E5", X"3A", X"48", X"5C", --1610
  X"E6", X"38", X"0F", X"0F", X"0F", X"F6", X"08", X"32", --1618
  X"90", X"6E", X"1A", X"13", X"B7", X"28", X"09", X"6F", --1620
  X"1A", X"13", X"67", X"CD", X"39", X"16", X"18", X"F2", --1628
  X"E1", X"F1", X"C1", X"D5", X"ED", X"5B", X"8E", X"6E", --1630
  X"C9", X"CD", X"40", X"16", X"2D", X"20", X"FA", X"C9", --1638
  X"3A", X"90", X"6E", X"CD", X"4A", X"16", X"06", X"04", --1640
  X"10", X"FE", X"44", X"00", X"00", X"00", X"10", X"FB", --1648
  X"EE", X"10", X"D3", X"FE", X"C9", X"00", X"01", X"02", --1650
  X"02", X"03", X"04", X"05", X"05", X"06", X"07", X"08", --1658
  X"09", X"09", X"0A", X"0B", X"0C", X"0C", X"0D", X"0E", --1660
  X"0F", X"10", X"10", X"11", X"12", X"13", X"13", X"14", --1668
  X"15", X"16", X"17", X"17", X"18", X"19", X"1A", X"1A", --1670
  X"1B", X"1C", X"1D", X"1D", X"1E", X"1F", X"20", X"20", --1678
  X"21", X"22", X"23", X"24", X"24", X"25", X"26", X"27", --1680
  X"27", X"28", X"29", X"29", X"2A", X"2B", X"2C", X"2C", --1688
  X"2D", X"2E", X"2F", X"2F", X"30", X"31", X"32", X"32", --1690
  X"33", X"34", X"34", X"35", X"36", X"36", X"37", X"38", --1698
  X"39", X"39", X"3A", X"3B", X"3B", X"3C", X"3D", X"3D", --16A0
  X"3E", X"3F", X"40", X"40", X"41", X"42", X"42", X"43", --16A8
  X"44", X"44", X"45", X"45", X"46", X"47", X"47", X"48", --16B0
  X"49", X"49", X"4A", X"4B", X"4B", X"4C", X"4D", X"4D", --16B8
  X"4E", X"4E", X"4F", X"50", X"50", X"51", X"51", X"52", --16C0
  X"53", X"53", X"54", X"54", X"55", X"56", X"56", X"57", --16C8
  X"57", X"58", X"58", X"59", X"5A", X"5A", X"5B", X"5B", --16D0
  X"5C", X"5C", X"5D", X"5D", X"5E", X"5E", X"5F", X"5F", --16D8
  X"60", X"60", X"61", X"61", X"62", X"62", X"63", X"63", --16E0
  X"64", X"64", X"65", X"65", X"66", X"66", X"67", X"67", --16E8
  X"68", X"68", X"69", X"69", X"69", X"6A", X"6A", X"6B", --16F0
  X"6B", X"6C", X"6C", X"6C", X"6D", X"6D", X"6E", X"6E", --16F8
  X"6E", X"6F", X"6F", X"70", X"70", X"70", X"71", X"71", --1700
  X"71", X"72", X"72", X"72", X"73", X"73", X"73", X"74", --1708
  X"74", X"74", X"75", X"75", X"75", X"76", X"76", X"76", --1710
  X"76", X"77", X"77", X"77", X"78", X"78", X"78", X"78", --1718
  X"79", X"79", X"79", X"79", X"79", X"7A", X"7A", X"7A", --1720
  X"7A", X"7B", X"7B", X"7B", X"7B", X"7B", X"7C", X"7C", --1728
  X"7C", X"7C", X"7C", X"7C", X"7D", X"7D", X"7D", X"7D", --1730
  X"7D", X"7D", X"7D", X"7D", X"7E", X"7E", X"7E", X"7E", --1738
  X"7E", X"7E", X"7E", X"7E", X"7E", X"7E", X"7F", X"7F", --1740
  X"7F", X"7F", X"7F", X"7F", X"7F", X"7F", X"7F", X"7F", --1748
  X"7F", X"7F", X"7F", X"7F", X"7F", X"01", X"FC", X"03", --1750
  X"CB", X"7C", X"28", X"04", X"09", X"30", X"FD", X"C9", --1758
  X"B7", X"ED", X"42", X"30", X"FC", X"09", X"C9", X"CD", --1760
  X"55", X"17", X"01", X"FF", X"00", X"B7", X"ED", X"42", --1768
  X"30", X"03", X"09", X"18", X"21", X"ED", X"42", X"30", --1770
  X"08", X"7D", X"ED", X"44", X"6F", X"26", X"00", X"18", --1778
  X"15", X"ED", X"42", X"38", X"0A", X"ED", X"42", X"7D", --1780
  X"ED", X"44", X"6F", X"26", X"00", X"18", X"01", X"09", --1788
  X"CD", X"96", X"17", X"ED", X"44", X"C9", X"01", X"55", --1790
  X"16", X"09", X"7E", X"C9", X"24", X"2B", X"C3", X"67", --1798
  X"17", X"2A", X"A2", X"6E", X"7E", X"23", X"22", X"91", --17A0
  X"6E", X"6F", X"3C", X"C8", X"26", X"00", X"29", X"29", --17A8
  X"29", X"ED", X"4B", X"1A", X"60", X"09", X"3E", X"08", --17B0
  X"32", X"95", X"6E", X"3A", X"9E", X"6E", X"32", X"9A", --17B8
  X"6E", X"3A", X"9D", X"6E", X"32", X"99", X"6E", X"3E", --17C0
  X"09", X"32", X"96", X"6E", X"7E", X"23", X"22", X"93", --17C8
  X"6E", X"07", X"32", X"97", X"6E", X"3A", X"96", X"6E", --17D0
  X"3D", X"20", X"32", X"3A", X"95", X"6E", X"3D", X"20", --17D8
  X"18", X"3A", X"A1", X"6E", X"47", X"3A", X"9F", X"6E", --17E0
  X"4F", X"3A", X"9D", X"6E", X"81", X"05", X"20", X"FC", --17E8
  X"32", X"9D", X"6E", X"2A", X"91", X"6E", X"C3", X"A4", --17F0
  X"17", X"32", X"95", X"6E", X"3A", X"A0", X"6E", X"47", --17F8
  X"3A", X"9A", X"6E", X"80", X"32", X"9A", X"6E", X"2A", --1800
  X"93", X"6E", X"C3", X"C1", X"17", X"32", X"96", X"6E", --1808
  X"3A", X"9F", X"6E", X"47", X"3A", X"9A", X"6E", X"32", --1810
  X"98", X"6E", X"3A", X"A0", X"6E", X"4F", X"C5", X"CD", --1818
  X"45", X"18", X"C1", X"3A", X"98", X"6E", X"3C", X"32", --1820
  X"98", X"6E", X"0D", X"20", X"F1", X"3A", X"99", X"6E", --1828
  X"3C", X"32", X"99", X"6E", X"05", X"20", X"DD", X"3A", --1830
  X"97", X"6E", X"C3", X"D1", X"17", X"80", X"40", X"20", --1838
  X"10", X"08", X"04", X"02", X"01", X"3A", X"9C", X"6E", --1840
  X"EE", X"FF", X"47", X"3A", X"9B", X"6E", X"A0", X"47", --1848
  X"3A", X"99", X"6E", X"E6", X"F8", X"6F", X"3A", X"98", --1850
  X"6E", X"FE", X"C0", X"D0", X"1F", X"1F", X"1F", X"E6", --1858
  X"1F", X"67", X"CB", X"1C", X"CB", X"1D", X"CB", X"1C", --1860
  X"CB", X"1D", X"CB", X"1C", X"CB", X"1D", X"3E", X"58", --1868
  X"B4", X"67", X"3A", X"9C", X"6E", X"A6", X"B0", X"77", --1870
  X"3A", X"98", X"6E", X"47", X"E6", X"07", X"F6", X"40", --1878
  X"67", X"78", X"1F", X"1F", X"1F", X"E6", X"18", X"B4", --1880
  X"67", X"78", X"17", X"17", X"E6", X"E0", X"6F", X"3A", --1888
  X"99", X"6E", X"47", X"1F", X"1F", X"1F", X"E6", X"1F", --1890
  X"B5", X"6F", X"EB", X"21", X"3D", X"18", X"78", X"E6", --1898
  X"07", X"4F", X"06", X"00", X"09", X"46", X"1A", X"21", --18A0
  X"97", X"6E", X"CB", X"46", X"28", X"03", X"B0", X"12", --18A8
  X"C9", X"2F", X"B0", X"2F", X"12", X"C9", X"2A", X"A6", --18B0
  X"6E", X"CB", X"15", X"CB", X"14", X"CB", X"15", X"CB", --18B8
  X"14", X"4C", X"3A", X"A4", X"6E", X"17", X"47", X"ED", --18C0
  X"5B", X"A5", X"6E", X"CB", X"13", X"CB", X"12", X"CB", --18C8
  X"BA", X"2A", X"A4", X"6E", X"09", X"22", X"A4", X"6E", --18D0
  X"2A", X"A6", X"6E", X"ED", X"5A", X"CB", X"BC", X"22", --18D8
  X"A6", X"6E", X"F0", X"21", X"A4", X"6E", X"34", X"C0", --18E0
  X"34", X"18", X"FB", X"C5", X"6F", X"26", X"00", X"29", --18E8
  X"29", X"29", X"ED", X"4B", X"1A", X"60", X"09", X"C1", --18F0
  X"C9", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --18F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1900
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1908
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1910
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1918
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1920
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1928
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1930
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1938
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1940
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1948
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1950
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1958
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1960
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1968
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1970
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1978
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1980
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1988
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1990
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1998
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --19A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --19A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --19B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --19B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --19C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --19C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --19D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --19D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --19E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --19E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --19F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --19F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1A98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1AA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1AA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1AB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1AB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1AC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1AC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1AD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1AD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1AE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1AE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1AF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1AF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1B98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1BA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1BA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1BB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1BB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1BC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1BC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1BD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1BD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1BE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1BE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1BF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1BF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1C98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1CA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1CA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1CB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1CB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1CC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1CC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1CD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1CD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1CE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1CE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1CF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1CF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1D98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1DA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1DA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1DB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1DB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1DC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1DC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1DD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1DD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1DE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1DE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1DF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1DF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1E98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1EA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1EA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1EB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1EB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1EC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1EC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1ED0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1ED8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1EE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1EE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1EF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1EF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1F98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1FA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1FA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1FB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1FB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1FC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1FC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1FD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1FD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1FE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1FE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1FF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1FF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2000
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2008
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2010
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2018
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2020
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2028
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2030
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2038
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2040
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2048
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2050
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2058
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2060
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2068
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2070
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2078
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2080
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2088
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2090
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2098
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --20A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --20A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --20B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --20B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --20C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --20C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --20D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --20D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --20E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --20E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --20F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --20F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2100
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2108
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2110
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2118
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2120
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2128
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2130
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2138
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2140
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2148
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2150
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2158
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2160
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2168
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2170
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2178
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2180
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2188
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2190
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2198
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --21A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --21A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --21B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --21B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --21C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --21C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --21D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --21D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --21E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --21E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --21F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --21F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2200
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2208
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2210
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2218
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2220
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2228
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2230
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2238
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2240
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2248
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2250
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2258
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2260
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2268
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2270
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2278
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2280
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2288
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2290
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2298
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --22A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --22A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --22B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --22B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --22C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --22C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --22D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --22D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --22E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --22E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --22F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --22F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2300
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2308
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2310
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2318
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2320
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2328
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2330
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2338
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2340
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2348
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2350
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2358
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2360
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2368
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2370
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2378
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2380
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2388
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2390
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2398
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --23A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --23A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --23B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --23B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --23C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --23C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --23D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --23D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --23E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --23E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --23F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --23F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2400
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2408
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2410
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2418
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2420
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2428
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2430
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2438
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2440
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2448
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2450
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2458
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2460
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2468
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2470
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2478
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2480
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2488
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2490
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2498
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --24A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --24A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --24B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --24B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --24C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --24C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --24D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --24D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --24E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --24E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --24F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --24F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2500
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2508
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2510
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2518
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2520
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2528
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2530
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2538
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2540
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2548
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2550
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2558
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2560
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2568
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2570
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2578
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2580
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2588
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2590
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2598
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --25A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --25A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --25B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --25B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --25C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --25C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --25D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --25D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --25E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --25E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --25F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --25F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2600
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2608
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2610
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2618
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2620
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2628
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2630
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2638
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2640
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2648
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2650
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2658
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2660
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2668
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2670
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2678
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2680
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2688
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2690
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2698
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --26A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --26A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --26B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --26B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --26C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --26C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --26D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --26D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --26E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --26E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --26F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --26F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2700
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2708
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2710
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2718
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2720
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2728
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2730
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2738
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2740
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2748
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2750
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2758
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2760
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2768
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2770
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2778
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2780
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2788
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2790
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2798
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --27A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --27A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --27B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --27B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --27C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --27C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --27D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --27D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --27E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --27E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --27F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --27F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2800
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2808
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2810
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2818
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2820
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2828
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2830
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2838
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2840
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2848
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2850
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2858
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2860
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2868
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2870
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2878
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2880
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2888
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2890
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2898
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --28A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --28A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --28B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --28B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --28C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --28C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --28D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --28D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --28E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --28E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --28F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --28F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2900
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2908
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2910
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2918
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2920
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2928
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2930
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2938
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2940
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2948
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2950
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2958
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2960
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2968
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2970
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2978
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2980
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2988
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2990
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2998
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --29A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --29A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --29B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --29B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --29C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --29C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --29D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --29D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --29E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --29E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --29F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --29F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2A98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2AA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2AA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2AB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2AB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2AC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2AC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2AD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2AD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2AE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2AE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2AF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2AF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2B98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2BA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2BA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2BB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2BB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2BC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2BC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2BD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2BD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2BE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2BE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2BF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2BF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2C98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2CA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2CA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2CB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2CB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2CC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2CC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2CD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2CD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2CE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2CE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2CF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2CF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2D98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2DA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2DA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2DB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2DB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2DC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2DC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2DD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2DD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2DE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2DE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2DF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2DF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2E98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2EA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2EA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2EB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2EB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2EC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2EC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2ED0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2ED8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2EE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2EE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2EF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2EF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2F98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2FA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2FA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2FB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2FB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2FC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2FC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2FD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2FD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2FE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2FE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2FF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --2FF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3000
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3008
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3010
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3018
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3020
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3028
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3030
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3038
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3040
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3048
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3050
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3058
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3060
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3068
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3070
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3078
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3080
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3088
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3090
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3098
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --30A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --30A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --30B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --30B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --30C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --30C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --30D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --30D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --30E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --30E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --30F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --30F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3100
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3108
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3110
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3118
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3120
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3128
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3130
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3138
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3140
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3148
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3150
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3158
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3160
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3168
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3170
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3178
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3180
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3188
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3190
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3198
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --31A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --31A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --31B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --31B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --31C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --31C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --31D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --31D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --31E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --31E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --31F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --31F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3200
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3208
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3210
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3218
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3220
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3228
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3230
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3238
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3240
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3248
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3250
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3258
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3260
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3268
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3270
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3278
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3280
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3288
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3290
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3298
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --32A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --32A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --32B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --32B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --32C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --32C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --32D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --32D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --32E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --32E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --32F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --32F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3300
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3308
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3310
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3318
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3320
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3328
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3330
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3338
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3340
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3348
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3350
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3358
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3360
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3368
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3370
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3378
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3380
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3388
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3390
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3398
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --33A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --33A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --33B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --33B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --33C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --33C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --33D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --33D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --33E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --33E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --33F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --33F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3400
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3408
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3410
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3418
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3420
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3428
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3430
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3438
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3440
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3448
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3450
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3458
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3460
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3468
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3470
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3478
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3480
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3488
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3490
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3498
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --34A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --34A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --34B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --34B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --34C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --34C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --34D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --34D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --34E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --34E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --34F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --34F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3500
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3508
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3510
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3518
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3520
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3528
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3530
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3538
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3540
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3548
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3550
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3558
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3560
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3568
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3570
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3578
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3580
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3588
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3590
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3598
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --35A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --35A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --35B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --35B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --35C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --35C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --35D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --35D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --35E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --35E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --35F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --35F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3600
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3608
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3610
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3618
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3620
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3628
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3630
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3638
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3640
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3648
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3650
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3658
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3660
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3668
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3670
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3678
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3680
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3688
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3690
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3698
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --36A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --36A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --36B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --36B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --36C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --36C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --36D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --36D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --36E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --36E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --36F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --36F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3700
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3708
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3710
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3718
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3720
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3728
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3730
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3738
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3740
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3748
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3750
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3758
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3760
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3768
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3770
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3778
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3780
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3788
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3790
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3798
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --37A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --37A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --37B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --37B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --37C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --37C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --37D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --37D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --37E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --37E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --37F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --37F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3800
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3808
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3810
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3818
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3820
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3828
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3830
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3838
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3840
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3848
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3850
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3858
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3860
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3868
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3870
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3878
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3880
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3888
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3890
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3898
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3900
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3908
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3910
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3918
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3920
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3928
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3930
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3938
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3940
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3948
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3950
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3958
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3960
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3968
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3970
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3978
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3980
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3988
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3990
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3998
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3D98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3DA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3DA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3DB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3DB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3DC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3DC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3DD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3DD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3DE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3DE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3DF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3DF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3E98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3EA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3EA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3EB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3EB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3EC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3EC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3ED0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3ED8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3EE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3EE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3EF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3EF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3F98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3FA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3FA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3FB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3FB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3FC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3FC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3FD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3FD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3FE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3FE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3FF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF");--3FF8

begin

  process (clk)
  begin
    if rising_edge(clk) then
      dout <= rom(to_integer(unsigned(addr)));
    end if;
  end process;

end architecture;
