library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

entity rom is port(
    clk     : in  std_logic;
    en      : in  std_logic;
    addr    : in  std_logic_vector(13 downto 0);
    dataout : out std_logic_vector( 7 downto 0));
end vram;

architecture Behavioral of vram is

  type arrena is array(7 downto 0) of std_logic;
  type arrdoa is array(7 downto 0) of std_logic_vector(7 downto 0);
  signal ena : arrena;
  signal doa : arrdoa;

begin
  process(addr, en, doa)
  variable i : integer;
  begin
    dataout <= (others => '0');
    for i in 0 to 7 loop
      ena(i) <= '0';
      if en='1' and to_integer(unsigned(addr(12 downto 11))) = i then
        ena(i) <= '1';
        dataout <= doa(i);
      end if;
    end loop;
  end process;

  rom0 : RAMB16_S9
  generic map (
    init_00 => X"D0007DCD7E5C5D2AFFFFFFFFFF15F2C343185C5F225C5D2A11CBC3FFFF11AFF3",
    init_01 => X"7822235C782AE5F5169EC3E55C612AC5FFFFFFFFFF335BC3FFFFFFF7180074CD",
    init_02 => X"FF16C5C35C3D7BED0075FD6EE1C9FBF1E1C1D102BFCDD5C54034FD0320B57C5C",
    init_03 => X"D021FEC97E5C5D22235C5D2A45EDF1E1E90120B57C5CB02AE5F5FFFFFFFFFFFF",
    init_04 => X"50A459454B4E49C44E52BFC95C5D223723013816FE23D83F18FED810FEC80DFE",
    init_05 => X"C5444F43A44C4156C24154D441D2545441A44E4545524353D44E494F50CE46C9",
    init_06 => X"D44E49D05845CE4CCE5441D34341CE5341CE4154D34F43CE4953CE454CCC4156",
    init_07 => X"CE4942D44F4EA4524843A4525453D25355CE49CB454550D34241CE4753D25153",
    init_08 => X"43CE4620464544D0455453CF54CE454854C54E494CBE3CBD3EBD3CC44E41D24F",
    init_09 => X"454DA32045534F4C43A3204E45504FC553415245C5564F4DD4414D524F46D441",
    init_0A => X"C853414C46D245504150CB4E49C54C43524943D0454542D94649524556C54752",
    init_0B => X"53D453494C4CD44E4952504CD4554FD245564FC5535245564E49D44847495242",
    init_0C => X"49544E4F43D24544524F42D7454EC5524F54534552C1544144C4414552D04F54",
    init_0D => X"C4414F4CD455504E49C25553204F47CF54204F47D24F46CD4552CD4944C5554E",
    init_0E => X"CE5552D44F4C50D44E495250C54B4F50D458454EC553554150D4454CD453494C",
    init_0F => X"5255544552D241454C43D7415244D34C43C649C55A494D4F444E4152C5564153",
    init_10 => X"4F4C0E5844453338494B4D4346523437554A4E5647543536594842D9504F43CE",
    init_11 => X"A5E5BAB2ADBEA6A7C0B1B0AFBBBDBCB4E4E0C4E341513130500D205A53573239",
    init_12 => X"D75BD9B6DB5DD57CD6B57FDFDEDDABAAAEBFD87D7BB75CDADC7EB8C1B9B3E1C2",
    init_13 => X"2FC53EC33CC7223B2C2E3D2B2DAC5ECBCCC8CD3F2AE20F090B0A08050406070C",
    init_14 => X"147D670E281FE62F78EDFEFE01FFFF112F2ECFA9D2D1D4D3CAA8CED03AC660C9",
    init_15 => X"CDC918FE575A7BC819FEC828FEC83C7AE63800CB2DF4205F53FA303CCB08D6C0",
    init_16 => X"BE5C0021D0031ECDEE20BD5C04217DFF3602202B352307207ECB5C0021C0028E",
    init_17 => X"FD074EFD23775C093A23053623775FC87ECBEB04207ECB2728BE5C0421EB2E28",
    init_18 => X"1642EA187E23775C0A3AC03523053623C9EE01CBFD5C083277E10333CDE50156",
    init_19 => X"4FC60328034FFA0D2F383AFE7BC9377E19020521C078CB032018FED027FE7B00",
    init_1A => X"04C05E30CBFD0A285ACBF42840CB022921C97E19001602052103280401EB21C9",
    init_1B => X"C6C80420D6073038FED32868CB0254211920039DFA0DD830FEC9A5C6C920C6C0",
    init_1C => X"CBC804C90FEEC80480C607E6B62830FEBA2839FE023021C9FEC6C80436D6C908",
    init_1D => X"064F03E62F3DCB3DCB7DF3C9403EC95F3EC020FE062822FE10D6A42002302168",
    init_1E => X"EE03D6C2053F0EFD200D0C0400000008F60F0F0F38E65C483A09DD03D121DD00",
    init_1F => X"6CEC3403C02731EFC9FBE9DD0C4DE9DD1B4D790928B37A092067CB4F44FED310",
    init_20 => X"F23CC6785020BE235420B99F177846234E235E20A77E5C9221380FA104F51F98",
    init_21 => X"C0EF7786F13804EF33B4CD3406CD046E21C50CC6FB300CD604FA06046CE20425",
    init_22 => X"CDC51E99CD38037135340501809F55438034E004E0EF22300BFE1E94CD383102",
    init_23 => X"901B891F17D512897560970A898612D002890ACF03B5C31BC8B37A5950E11E99",
    init_24 => X"0000005C895400A74F89736AFF43893E49FF3889B1369D2E89CA53D024890241",
    init_25 => X"CB09F80D6B622BF1CDE5D0E11C8AFA875C3B3A24FBCD0510F1768924F6146989",
    init_26 => X"A4060FEEFED3FE1047023EF32BDD13080C982103287FCB1F8021E5053F21C9FE",
    init_27 => X"B37A0507C36F083B0E01FED3FE1037060D3EFED3FE102F0604D8F22505F5202D",
    init_28 => X"3E06FED3FE1042060430FE1078CB79F4186C0525C337013E67AD7C006EDD0C28",
    init_29 => X"F5C9FE103B0604FEC23C7AD01FFEDB7F3E310623DD1B0514C215CB3CAF05EF20",
    init_2A => X"3F21FED30F3EF3150814C9F10CCF0238FB1FFEDB7F3EFED30F0F0F38E65C483A",
    init_2B => X"EB3005E3CDF920B57C2BFE10041521FA3005E7CDC0BF4F02F620E61FFEDBE505",
    init_2C => X"79D005E7CDF430D4FE78D53005E7CDC906F12024E030B8C63EE43005E3CD9C06",
    init_2D => X"007EDD0718134F1F79C0AD11CB0F180075DD0F300720081F18B00600264F03EE",
    init_2E => X"7CCA20B37A67AD7C05CAD2B00615CBB8CB3ED005E3CD012EB206081B23DDC0AD",
    init_2F => X"F607E64F2F79F32820E6A9D01FFEDB7F3EC804A7FD203D163ED005E7CDC901FE",
    init_30 => X"0E0228A75C743A0011013C282530CD1C8CCD5C7432E0D65C743AF1C937FED308",
    init_31 => X"A75C743A0F3003090BFFF6212BF1CDFF0136DDFC101312203E0B06E1DDD5F722",
    init_32 => X"E71C8ACA03FE5C743A4920E4FEDFB0EDEB23E1E5DD000A010A28B1780ECF0220",
    init_33 => X"230B77DD7E2318282530CD1C8AC201CF15283D5C743A0000210B30F9CB28B2CD",
    init_34 => X"075AC3EB1BEECDE7DA2029FEE7EB0077DD3C012871CB013E0E71DD230C77DD7E",
    init_35 => X"74DD0D75DD4000211B0C36DD000B36DD1BEECDE71C8ACA03FE5C743A1F20AAFE",
    init_36 => X"181CE6CD1C8ACAA75C743A0C202048CDE71C8ACA03FE5C743A4F20AFFE4D180E",
    init_37 => X"DD1E99CD1BEECD1C82CDE704181CE6CD1C8ACAA75C743A0C282CFEDF1C82CD0F",
    init_38 => X"0E36DD1BEECD0928CAFE4418030036DD69600E70DD0D71DD1E99CD0C70DD0B71",
    init_39 => X"592A000036DD0E70DD0D71DD1E99CD1BEECD1C82CDE71C8AC2A75C743A171880",
    init_3A => X"70CAA75C743AEB1074DD0F75DD52ED5C4B2A0C74DD0B75DD52ED375C535BED5C",
    init_3B => X"800E035236FD1601CDFE3EF230E1DD0556CD37AF001111E5DD09DD001101E509",
    init_3C => X"7E0A0619FFF021D1E5DDC10C0ACDC509C011D93004FEF60E0220EFBEDD007EDD",
    init_3D => X"3A0C2803FE007EDDE1D70D3EB32079CBF610D70C012023BE1A134F807903203C",
    init_3E => X"263852ED0D28B57C0C56DD0B5EDDFB66DDFA6EDDE508B6CA02FE0808CA3D5C74",
    init_3F => X"A701203702FE5C743AE1DDE50E66DD0D6EDD0620B57CE11D2003FE007EDD0728",
    write_mode => "READ_FIRST")
  port map (
    do    => doa(0),
    addr  => addr(10 downto 0),
    clk   => clk,
    en    => ena(0),
    we    => '0',
    ssr   => '0');

  rom1 : RAMB16_S9
  generic map (
    init_00 => X"EBFB66DDFA6EDD0C18EB1313130620B57CE50C56DD0B5EDD1ACFD80556CDFF3E",
    init_01 => X"03032B4E2B462B1328B57C3E28A7007EDDE11F05CD4D4419000511093852ED37",
    init_02 => X"55CDF5FD7EDD030303C50C46DD0B4EDD2B5C592A5C5F2ADD19E8CD5C5F22DD03",
    init_03 => X"DD0B4EDD5C5F22DD2B5C592AEB0802C3FF3E37E1DDE52372237323D177F12316",
    init_04 => X"E67C0E66DD5C4B22091046DD0F4EDD235C5F2ADD1655CDC5E5C119E5CDC50C46",
    init_05 => X"36F703C50C46DD0B4EDD0802C3FF3E37E1DDD1000A36FD5C42220D6EDD0A20C0",
    init_06 => X"1BBE1A022023BE131A1920C0E67E5C535BEDE10802CDFF3E37E1DDE5E5D1EB80",
    init_07 => X"28B9252880FE7E5C4B2AE5C880FE4F7EE218092CCDEC18E119B8CDEBE508302B",
    init_08 => X"18E10318E1F730170620BE1A1323E5D5D11220A0FEE0E6F018EBC119B8CDC508",
    init_09 => X"D508085C5F2AEB19E8CD19B8CDEB5C5F22081020C418092CCD373CEBD1FF3EE0",
    init_0A => X"ED5C5353EDD1C1231655CD0318231655CD2B073808C5E35C532A5C5F2219B8CD",
    init_0B => X"02CBFD0C0ACD09A111AF1601CDFD3EE5C9D119E8CDD5C1E1B0EDEBD5C55C5F5B",
    init_0C => X"C2C3E1DDFF3E0C56DD0B5EDDFD10763206E1DD04C2CDAF001111E5DD15D4CDEE",
    init_0D => X"79656B20796E61207373657270206E656874202C657061742074726174538004",
    init_0E => X"61726168430DA03A7961727261207265626D754E0DA03A6D6172676F72500DAE",
    init_0F => X"693806FE0AD9D220FE0B03CDA03A73657479420DA03A79617272612072657463",
    init_10 => X"5B5C5D5E5F4F50375253542910574E0B03C3E5195E1900165F0A0B21653018FE",
    init_11 => X"5C913A0DD9C3210E050320B8183E020E0409204E01CBFD1120B9223E0C53545A",
    init_12 => X"CD0DD9C3050C55CD210E0ECDC24E01CBFDC95C9132F10B65CD203E015736FDF5",
    init_13 => X"5C0E320A871103180A6D110B185C0F320A87116C183F3E5A1810E63D3D790B03",
    init_14 => X"0C38911F3E4A4429202211DA16FE7D575C0E2A0A80CD09F411C97223735C512A",
    init_15 => X"C30C86DA31BEFD0C55C24602CBFD04473C1E9FDA90163E16204E01CBFD4F02C6",
    init_16 => X"4E01CBFD0B24CDC9F820150C3BCD203EC601CBFD57C81FE63D810B03CD7C0DD9",
    init_17 => X"224571FDC95C86225C8243ED5C8A43EDC95C84225C8843ED08204602CBFD1A20",
    init_18 => X"454EFDC95C862A5C8A4BEDC84602CBFD5C842A5C884BED14204E01CBFDC95C80",
    init_19 => X"18CB0B3ECD5C922147185C92110B03CD0B38CD47263090FE3D3880FEC95C802A",
    init_1A => X"CD0B185C7B4BEDC515C60930A5D6C9FB200D2377040EB1F0E69F18CB4F0FE69F",
    init_1B => X"79EBC1092929296F0026C6CB022020FE86CB5C3B21EB5C364BEDC50B03C30C10",
    init_1C => X"FF065C913AE5C5D10C55CCD5B979D10ECDCDD506284E01CBFD4F050E20213E3D",
    init_1D => X"13380812A9AEA01A08EB37CE30CBFD05284E01CBFDA7083E4F9F1F1F0401381F",
    init_1E => X"E60F0F0F7CE618085F83203E08C9230DC1E10BDBCC4E01CBFD25EBF2203D2314",
    init_1F => X"08286657CBFD38EE022057CBC7E608287657CBFDABA2AB7E5C8F5BED6758F603",
    init_20 => X"CC4601CBFD203E09380C41CDF50095110418E30026E5C97707EE02206FCBF8E6",
    init_21 => X"D1D9D7D9D5203ED803FE7AD882FE032848FED1F53087131A0C3BCD7FE61A0C3B",
    init_22 => X"FD78D50DD911C04E01CBFDC941D61AD820FEF1EBF8203DFB28237ECB3CEBF5C9",
    init_23 => X"3F7BED1601CD003E5A281D2D5EFD16286602CBFDC01B3831BEFD0D02C24602CB",
    init_24 => X"1601CDFD3EF55C913AE55C8F2A5C8C3290183E45205235FD04CFC9A602CBFD5C",
    init_25 => X"F64128E2FE452820FED915D4CDD9AECBDECB5C3B21EE02CBFD0C0ACD0CF811AF",
    init_26 => X"7C0E9BCDC5210E043146FD0DFECD5C8F22E15C9132F11601CDFE3E3B286EFE20",
    init_27 => X"BF6C6C6F72637380C9C1FA1023137112EB20064E1A5AE0116758F603E60F0F0F",
    init_28 => X"5C6B21F5780D4DCDE55C912AE55C8F2A47C544EDD019D63186FD803802FE0CCF",
    init_29 => X"5C884BED5C8F22E15775FDE1E8203DF10E00CD1806340338BE5C8921773C7846",
    init_2A => X"91215C8F220E6EFD6704284602CBFD5C8D2AAFC9C1C602CBFD0DD9CD8602CBFD",
    init_2B => X"C0210E44CD3146FD0D4DCDC6CBAECB5C3C210DAFCDC977AE55E6AE0F7E02205C",
    init_2C => X"A709F4115C512A1601CDFD3E023136FDF710FB200D772B200E0718055C8D3A5A",
    init_2D => X"01CDFE3E0D94CD8630CBFD5C7D220000212A18172101F6383F10A81123722373",
    init_2E => X"4E01CBFD5B0021182101015236FD72237309F4115C512A0E44CD18060D4DCD16",
    init_2F => X"17060ADCC31900165F91213EC10E9BCD47C518D63186FD05284602CBFD781220",
    init_30 => X"47EB19FFE021EBB0ED3D002001EB19F8E021EB0C207807E678E5C5080E0E9BCD",
    init_31 => X"EB19FFE0210E88CDCD200DC124E1DB20F8E6090706B0ED0006784F0F0F0F07E6",
    init_32 => X"0111B0ED1300365D540D0006784F0F0F0F07E678E5C5080E0E9BCDC50106B0ED",
    init_33 => X"5C483A03284602CBFD5C8D3A136B620E88CDDC200DC124E1E52047F8E63D1907",
    init_34 => X"0F5790183EC94D4429292929296861EB6750F63D0F0F0F7CC9210EC1B0ED0B77",
    init_35 => X"7D0A2007E67C24E1C10EF4CDC5E5400021B006F3C96740F618E67A6FE0E60F0F",
    init_36 => X"21FBFBD3043EF910C10EF4CDC508065B0021F30D18E7106784F8E69F3F6F20C6",
    init_37 => X"1F54CD57FBD302E69F03FE780DD9C3210E8E30CBFDFC10237747AF4675FD5B00",
    init_38 => X"FBDB1ACB13CB12CB0806235E200EEB30F887FBDB0CCF0EDFCDFBFBD3043E0A38",
    init_39 => X"5EFD0016F515D4CD5C3D73EDE5107F21E55C3D2AC9E9200DF010FBD37AFB301F",
    init_3A => X"0C3816FE570002013A3810FE2D3807FE313018FEE50F3821F103B5CD00C821FF",
    init_3B => X"1871237023C11655CD8607CBFD5C5B2AD515D4CD5F15D4CD101ECA7E37CBFD03",
    init_3C => X"C95C5B2AE5195E190F992100165FC95C5B53ED13121652CD5C5B2A8607CBFD0A",
    init_3D => X"23E51097CAB37A1695CD196ECD1097C26E37CBFD5C492AD4CF7E70B5506A6609",
    init_3E => X"55CD0F35FD2BE11601CDFF3EE5E35C512A1097CD1F05CD4D4409000A2146234E",
    init_3F => X"18190FCD5C492108206E37CBFDC91615CDE15C5B22232323235C592A0F34FD18",
    write_mode => "READ_FIRST")
  port map (
    do    => doa(1),
    addr  => addr(10 downto 0),
    clk   => clk,
    en    => ena(1),
    we    => '0',
    ssr   => '0');

  rom2 : RAMB16_S9
  generic map (
    init_00 => X"D4CD19E8C30001011031CDC95C5B2223C80DFE7E05181031CD1D18100036FD6D",
    init_01 => X"6B624D44C5D8C1231952ED1195CD37C9F9C07E00CBFD5C3D22E1E1E115D4CD15",
    init_02 => X"492AC06E37CBFDC9E638EB0942EDA723012000CE17D61A23092010FEF0E61A23",
    init_03 => X"FD0F81C3A8287E37CBFD1601C3003E1795CD191CCD5C4A211695CDEB196ECD5C",
    init_04 => X"2219E5CD2B1190CDE50F30C303B5CD1A9021FE5EFD0016FF0036FDA1286630CB",
    init_05 => X"02CBFDF5AE01CBFD5C083AC86E01CBFDA7111DC45E02CBFDC9E1000736FD5C5B",
    init_06 => X"5C6A2109202A1812C61F784F01E6470A3006FE2D3010FE523020FEF10D6EC46E",
    init_07 => X"103E4F07E647C9BFDE02CBFD0036022077BE5C41210DD6D80EFE0E1877AE083E",
    init_08 => X"0D4DCDC93772237323235C4F2A10A8115C0D3A0618110D11D371FD3C012058CB",
    init_09 => X"1195CD37E55C822A5C3D73EDE5116721E55C3D2AE55C8A2AAE02CBFD9E02CBFD",
    init_0A => X"203E1E305096FD7B06202638925C8B3A0D4DCDEBE35C8A2A18E1CDEB187DCDEB",
    init_0B => X"22E1E1D102185C8A5BEDFF0036FD03B5CD1A9021FE5EFD0016E918D109F4CDD5",
    init_0C => X"5BEDC86E37CBFD5C595BEDA72B5C612AC9002636FD5C8222E10DD9CDD5C15C3D",
    init_0D => X"EDD95CB25BEDFF3EF3C9F1200DFE237E19E8CC0006010EFE7EC95C632AD85C61",
    init_0E => X"BC2B02366B6200000000000047ED3F3EFED3073E47D95C7B2A5C385BED5CB44B",
    init_0F => X"192804D95C7B225C3853ED5CB443EDD92BF328350328350630231952EDA7FA20",
    init_10 => X"223C00215CB2225C3843ED0040012B5C7B2223EBB8EDEB00A8013EAF115CB422",
    init_11 => X"150115AF115C4F225CB621FB5C3A21FD56ED5C3D222B2BF92B3E365CB22A5C36",
    init_12 => X"225C6122238036230D365C59222380365C4B225C5322235C57222BEBB0EDEB00",
    init_13 => X"1115C621CA35FDC635FD5C09220523215C48325C8F325C8D32383E5C65225C63",
    init_14 => X"EE02CBFD0C0ACD153811AF0D6BCD023136FD0EDFCDCE01CBFDB0ED000E015C10",
    init_15 => X"30CBFD12207E00CBFD1B17CD0F2CCD1601CD003E16B0CD1795CD023136FD0718",
    init_16 => X"0DFEDF155DC2B17819FBCD5C5D225C592ADD18FF0036FD11A7CD5C592A402866",
    init_17 => X"010A36FDFF0036FDFE01CBFD5C8C324F96FD193E0D6ECD0DAFC44630CBFDC028",
    init_18 => X"5C0B222674FD3774FD000021F53C5C3A3A0ECDC44E30CBFDAE01CBFD761B8ACD",
    init_19 => X"3E15EFCD07C602380AFE47F1EE02CBFD0D6ECDAE37CBFD16B0CD5C1622000121",
    init_1A => X"CD00060D4EFDD73A3E1A1BCD5C454BED0C0ACD153611AF0C0ACD13911178D720",
    init_1B => X"CB5C44215C70110003010D34FD032015FE042809FE1B283C5C3A3A1097CD1A1B",
    init_1C => X"74756F68746977205458454ECB4F8012ACC39E01CBFDFF0A36FDB8ED0901287E",
    init_1D => X"20747069726373627553E46E756F6620746F6E20656C626169726156D24F4620",
    init_1E => X"4EEE656572637320666F2074754FF9726F6D656D20666F2074754FE76E6F7277",
    init_1F => X"55534F472074756F68746977204E5255544552E76962206F6F74207265626D75",
    init_20 => X"696C61766E49F46E656D657461747320504F5453E56C696620666F20646E45C2",
    init_21 => X"6F4EE5676E617220666F2074756F2072656765746E49F46E656D756772612064",
    init_22 => X"6570657220544E4F43202D204B41455242C349534142206E692065736E65736E",
    init_23 => X"4EE56D616E20656C69662064696C61766E49C154414420666F2074754FF37461",
    init_24 => X"20524F46D455504E49206E6920504F5453E56E696C20726F66206D6F6F72206F",
    init_25 => X"6E49E56369766564204F2F492064696C61766E49D458454E2074756F68746977",
    init_26 => X"4152ED6172676F7270206F746E69204B41455242F2756F6C6F632064696C6176",
    init_27 => X"696C61766E49F4736F6C20746E656D6574617453E46F6F67206F6E20504F544D",
    init_28 => X"20726574656D61726150C645442074756F68746977204E46ED61657274732064",
    init_29 => X"2032383931207FA02CF26F72726520676E6964616F6C2065706154F26F727265",
    init_2A => X"4943ED1313C3000001103EE4744C206863726165736552207269616C636E6953",
    init_2B => X"3D79C119E8CD19B8CD0620196ECD6960E552ED375C612AE5155521EB5C5D2A5C",
    init_2C => X"2AB8ED2B2B5C612A13C5C15C5322E11655CDD55C535BED2B03030303C52828B0",
    init_2D => X"09F45215C40F815315C409F44B10A809F412A2C3F1722B732B712B70C1EB5C49",
    init_2E => X"E6CDDE02CBFD04206E02CBFD0010000600010001000B0006000112CF805015C4",
    init_2F => X"D9E1162CCDEB56235E5C512AE5D983301E081823235C512AE5D907CFFA28D815",
    init_30 => X"23232323A630CBFD5C5122195C4F2A1B17CF0220B37A56235E5C266F16C687C9",
    init_31 => X"E630CBFDAE01CBFDC602CBFD001B501253064BE9195E0016D016DCCD162D214E",
    init_32 => X"5C652A1664CDE11F05CDE5000101C9CE01CBFD0D4DC38E01CBFD8602CBFD0418",
    init_33 => X"23D123732B72EB09EBD50930E31952EDA7E356235E0E3E5C4B21E5F5C9B8EDEB",
    init_34 => X"632AC95E2356F720C0E67E168F11EB0000C9EB19034D4452EDA7F1D1EBE8203D",
    init_35 => X"2A5C6122238036235C5B220D365C592AC923EBC15C6143EDC123231655CD2B5C",
    init_36 => X"B9C8A77E2319E5C35C595BEDC9E15C68225C9221E55C65225C632A5C63225C61",
    init_37 => X"702371EB46234E0915D401073819EBA3E2110000011701CD171ECDC937F82023",
    init_38 => X"94CDC9E101500353054BE90900064E16DCCD171621EB4E232323095C4F2AE5C9",
    init_39 => X"1628B178171ECD3801EFC92B46234E0900064F5C10210703C617CF023810FE1E",
    init_3A => X"F1CDE5C9722373175DCDCF2050FE042853FE08284BFEEB7E232323095C4F2AEB",
    init_3B => X"0A500853064BE9C10900064EF13016DCCD177A214FDFE61AC50ECF0220B1782B",
    init_3C => X"0DAFCD100236FD5C3F73ED9018C9E157D520B1780B101E0218061E0618011E00",
    init_3D => X"D522381952EDA75C6C5BED5C492AC630CBFD8602CBFD0E44CD3146FDC602CBFD",
    init_3E => X"185C6C53ED2B5E2356EB0E3809C119B8CDC5C1196ECDE352EDEB02C011196ECD",
    init_3F => X"CD000236FD023E0218033EC9A602CBFD1833CDEB0128196ECD5C6C2A5C6C22ED",
    write_mode => "READ_FIRST")
  port map (
    do    => doa(2),
    addr  => addr(10 downto 0),
    clk   => clk,
    en    => ena(2),
    we    => '0',
    ssr   => '0');

  rom3 : RAMB16_S9
  generic map (
    init_00 => X"CD03181CE6CD08181C82CDE706202CFE04283BFEDF14382070CDDF1601C42530",
    init_01 => X"3AF6286602CBFDD71855CD011E196ECD5C492269673FE6781E99CD1BEECD1CDE",
    init_02 => X"05283E161980CD5C494BEDE018E1D1190FCD5C6C21D5E5C8ABEE204F96FD5C6B",
    init_03 => X"01CBFDD70528A77A8601CBFD2323231A28CDC5D0C140FE7E2D73FD13CB000011",
    init_04 => X"C1CD3F3E052052EDA75C5F2AD6CB02286E37CBFD96CB5C3B219630CBFDEBD5C6",
    init_05 => X"7E232323232323C00EFEC9D1E0181937CDEB06280DFE2318B6CD7EEB18E1CD18",
    init_06 => X"D95C8F22E15774FDE109F4CD0036D5565C91215C8F22FDCBBCCBE55C8F2AD9C9",
    init_07 => X"DECB0B2856CB4B3E9ECB5C3B21161843C6042807CB5C413AC052EDA75C5B2AC9",
    init_08 => X"6E37CBFDE11695CD196ECD23EBE556235EC9D118C1CDD5433E02285E30CBFD3C",
    init_09 => X"2C3821FE30302D1BCD15EFC3F1283D42EDFC383C09AF0D18F8A77BC9732B72C0",
    init_0A => X"3AF50A2022FE0E1814285630CBFD16206E37CBFD0E203AFE2428CBFE9601CBFD",
    init_0B => X"F418EB19B8CDC5D01980CDC15D545C532AE5C9D7D601CBFDF15C6A3204EE5C6A",
    init_0C => X"5C5D2218B6CD7E23C9A70420BBE7C815000E5C5D22232323C9B92B7E23C0B87E",
    init_0D => X"6FCB173840FE7EE5C93715E3200DFEDF2841CB0420CBFE04283AFE0D012022FE",
    init_0E => X"52EDA7D1092346234E23230618FB307E2317120E02300005013F19C7FA871428",
    init_0F => X"222B5C592AC9E1B0EDD519E1EB1664CD034F2F79472F78C519DDCDC9EB194D44",
    init_10 => X"78CBAFE5D516C5C31C8ADA09D8F02104382DA2CD2D3BCD5C65225C9221E75C5D",
    init_11 => X"2ACDF60E192ACDFF9C01192ACDFC1801201EEBE55E2356D50818FF1E69602020",
    init_12 => X"706E6C2E817F9898989898989895929193B4AFC4BFBCCBB1C9D1E115EFCD7D19",
    init_13 => X"670006023D015D15445C490D426D3A512D432B590F4477371F172B413F569448",
    init_14 => X"051FCD051DAB00041D030506CC063D041F23001CEE001EED00061CF005CB061E",
    init_15 => X"6B001EAC031E5F001E4F031E80000817F9051EA10311B7001BB2052C02052089",
    init_16 => X"0B17F5051FC9050EAC00238205091E42031E27051DED051F3A000622DC00090D",
    init_17 => X"000A2C061F6005229400061E7A00080707070707072320050903F800080B0B0B",
    init_18 => X"32AF19FBCDBE01CBFD1793001793000A1793000A2C0A1793000A16E500061736",
    init_19 => X"1B7621EB283AFE7A280DFE0006DF1C8AFA0D34FD16BFCDE701185C3A323D5C47",
    init_1A => X"FE4FC51B52015C7422237E5C742A0318094E091A48214F1C8ADACED679E74FE5",
    init_1B => X"0ACBFD14CF02381F54CDC9E71C8AC2B9DFC905DFE5094E0900061C01210C3020",
    init_1C => X"6ECD33185C443A1B5C595BED2B5C612A5C4522FFFE2114287CCB5C422A71207E",
    init_1D => X"FEAFC0A6C03E5C552AC82530CDC1FFCF0F2878C0E67E474320A719285C443A19",
    init_1E => X"15FF0A36FD001E575C5D22EB5C55222319EB56235E235C4553ED5E235600CE01",
    init_1F => X"8AC31B28CA3AFEBA280DFEDFC1C1C02530CD16CF0828198BCD141B28CA0D72FD",
    init_20 => X"CDC9C5EB46234E5C742AEB1BEECCC1BF1CDECDCF81B4718E7B0B67094B1D0F1C",
    init_21 => X"2BF1C42530CDAF0D207601CBFD2996CC01CF1820CE37CBFD0830003736FD28B2",
    init_22 => X"56FDF124FBCDF55C3B3AC91BEECD1C56CDC1C95C4D225C7243EDEB77B65C7121",
    init_23 => X"202CFE1C82CDE7A918F114203C9FF679F528B2CDC92AFFC27ACB242040E6AA01",
    init_24 => X"4DC48602CBFD7E01CBFDF418C87601CBFD24FBCD0BCFC07601CBFD24FBCDE709",
    init_25 => X"30CDC977AEAAE6AE077E5C91215C8D225C8F2A1BEECD21FCCD13D65C743AF10D",
    init_26 => X"0DFE0605C39F1821E2CDDFB657CBFD77F8F67E5C90210D4DCD8602CBFD132825",
    init_27 => X"1BB3DA34E9CDEB3802EF0A282530CDC108CFC938A0EFC82530CD9C203AFE0428",
    init_28 => X"2AFFCD3801E00102C0EF38A1EF1BEECD06181BEECD1C82CDE70920CDFE1B29C3",
    init_29 => X"2AB0ED0A0EEBE1380202EFE5231655CD0D0E06380709000601FECB7E2B5C6822",
    init_2A => X"2A5744ED5C473A5C42225C452A3846FDD01DDACD7223140D56FD722373EB5C45",
    init_2B => X"92013EE7E818E70328B820F6E71138C15C5543ED1D86CD5C554BEDC5F31E5C5D",
    init_2C => X"4D4409E546234E235C4243ED4E2346C037C0E67E2318283AFE7E11CFC95C4432",
    init_2D => X"E2E0EF5C6822231F287ECB5C4D2A1C2EC24E37CBFDE018D0C1198BCDC50016E1",
    init_2E => X"0036E2E0E1EF00CF1E73C3EB662356235E19000F115C682AD81DDACD3802C00F",
    init_2F => X"282CFE7E5C572A5C5F22DF29282530CD1C1FCDE7C93738C9A738040037030102",
    init_30 => X"FEDF0078CD002636FD5C5F2A5C5722DF1C56CD0077CD0DCF02301D86CDE41E09",
    init_31 => X"C3020011B9ED47E43EF518E71BEEC42CFE24FBCD0B202530CDC91BEECDC9282C",
    init_32 => X"2AC95C7643ED5C784BED0420B1781E99CDC95C57222B196ECD69601E99CD198B",
    init_33 => X"C979ED1E85CDC90A72FD5C42222C30F0FE7C001669601E99CD0C183656FD5C6E",
    init_34 => X"CFC801382DA2CD03182DD5CDC9F11E99CDF544ED022815382DD5CDC9021E85CD",
    init_35 => X"2B5C592A5C4B5BEDC55CB24BED0420B1781E99CD03181E45CD0000011E67CD0A",
    init_36 => X"5CB222EB15CF023052EDA75CB42A083052EDD1190032115C652A0D6BCD19E5CD",
    init_37 => X"CDD55C3D73EDE5C55C454BED33E3240D66FDD1E9EB5C3D73EDC5F92B3E36C1D1",
    init_38 => X"1F05CD0000010055C3032ED872ED033819005021EB0A38095C652A0014011E67",
    init_39 => X"780B761E99CD06CFE5D51E73C3C55C3D73EDEBE33B0B283EFE7AD1E1C1C94D44",
    init_3A => X"C91FFEDBFE3ED81FFEDB7F3EC9AE01CBFDEE286E01CBFD0301203CA1780C28B1",
    init_3B => X"2028FEE7B601CBFD052024FEE716302C8DCDF601CBFD1E39C3CE3E05282530CD",
    init_3C => X"FE0E3623231655CD000601EBE7EB022024FEE7EB1C8AD22C8DCD202829FEE73C",
    init_3D => X"1C8AC240E601AEFDF124FBCDF55C3B3AE70E203DFEE7132029FEE018E703202C",
    init_3E => X"DFC91BEECD1FDFCD0D4DCD1601C42530CD023E0218033EE9C8E12530CD1BEECD",
    init_3F => X"20ACFEDFC9D70D3E1FC3CDC829FEF328204ECD1FFCCDFB28204ECD0D282045CD",
    write_mode => "READ_FIRST")
  port map (
    do    => doa(3),
    addr  => addr(10 downto 0),
    clk   => clk,
    en    => ena(3),
    we    => '0',
    ssr   => '0');

  rom4 : RAMB16_S9
  generic map (
    init_00 => X"79D7173E1E99CD1FC3CD1C82CDE71220ADFE1018163E2307CD1FC3CD1C79CD0D",
    init_01 => X"C80BB1782DE3C22BF1CC7601CBFD1FC3CD24FBCDD02070CDD021F2CDC9D778D7",
    init_02 => X"18D7063E0B282530CD0A202CFE14283BFEDFC93AFEC80DFEC829FEF718D7131A",
    init_03 => X"FE1E94CD1FC3CDA71C82CDE7C03723FEC9BFC101202045CDE71FF5CDC027FE06",
    init_04 => X"1BEECD20C1CD010236FD0D6ECD1601CD013E08282530CDC9A71601CD160ED210",
    init_05 => X"6EC30DD9CD8602CBFD5C8C3290193E5C8843ED47210E0338B85C6B3A5C884BED",
    init_06 => X"1C1FCDE71120CAFE21B2C3E71C8AC229FEDF1FDFCDE70E2028FEFB28204ECD0D",
    init_07 => X"21B2CA2530CDBE37CBFD1C1FCD21AFD22C8DCD0D181C8AC27601CBFDFE37CBFD",
    init_08 => X"790D36F777B6030E022040E65C3B3A0B207ECB000101EECBB6CB5C712116BFCD",
    init_09 => X"CBFDE5213A21E55C3D2AE55C5D2A2C207E37CBFD5C5B22772B12223E05300F0F",
    init_0A => X"2CCD031821B9CDBE01CBFD0F2CCDFF0036FD11A7CD5C612A5C3D73ED04286630",
    init_0B => X"E11C20BECB7ECBAECB5C71210DD9CD5C824BED111DCD0A2021D6CD002236FD0F",
    init_0C => X"5BED5C632A17185C5D22002636FD5C5F2A21B9CDFE01CBFD5C5F22E15C3D22E1",
    init_0D => X"DF5C5D225C612AC920C1CA204ECD1FFCCD03182AFFCD2AB2CD4D4452ED375C61",
    init_0E => X"4BFE7E232323235C512A10CFC82530CD0BCFC80DFEDF1C59CD5C713A0C28E2FE",
    init_0F => X"CDF5C9D6F1E7F5D83FDFFED8D9FE1C8AC3F2283BFEF6282CFEDFD821F2CDE7C9",
    init_10 => X"7A01FE562800CE02D61D2800CE11D6C9D77AD7F1571E94CDF51FC3CDA7F11C82",
    init_11 => X"7A4F3806070707053807067A38185C912179163002FE7A4F0406070704200106",
    init_12 => X"9FBA073E226CCD794F78012824E62FB007287E0B3808FE5C8F2113CF02380AFE",
    init_13 => X"FE7A4F40060F032080060F7A9FC9782377AEA0AE9FBA083E4750E60707226CCD",
    init_14 => X"070707FED3A93008FE1E94CDD8180F0F0F79226CCD5C8F2179BD3002FE042808",
    init_15 => X"0707077967A8F8E6A81FA71F371FA74724F9DA90AF3EC95C483207EE02206FCB",
    init_16 => X"CD2307CD2D28C301E6FD10077E044722AACD2307CDC907E6796F0707A8C7E6A8",
    init_17 => X"2051CBA0012041CB574EFD7E47FD100FFE3E044722AACD5C7D43ED0D4DC322E5",
    init_18 => X"C9FF0EC8010E24F9DA2DD5CDC94F51C1592314CDC5472314CD0BDBC3772FA802",
    init_19 => X"833638A3EFA1183802EF053081FE7E383D2AEF1BEECD1C82CDE71C8AC22CFEDF",
    init_1A => X"0302C001C2EF22DCC3C1380202EF083080FE7E3804E131EFC5247DCD3802C5EF",
    init_1B => X"C3C15C7D2267E11E94CDE56F1E94CD6234FD3802C1A0E03101E03101C00FE001",
    init_1C => X"380206003030311F04A2C5EF1BEECD1C82CDE72477C31BEECD06282CFEDF2420",
    init_1D => X"77C3380202EF073081FE7E383D01E02A05E00F2AE101E12A3102C102C02477C3",
    init_1E => X"02C51F3104A203E0E5E204E1310102C204E1310102C10501E102EFC5247DCD24",
    init_1F => X"81FE1A38020F2AE12AC20304E5E204E002C101E10F04E2E004E5C102C202C020",
    init_20 => X"C138E5E00FC5EF2D28CD5C7E3A38010FC0EF2D28CD5C7D3A3801EFC52477DAC1",
    init_21 => X"310FE102C0EFC53802C20F04E3E204E402C10304E4E204E331E1EF14183C2805",
    init_22 => X"EFC610C124B7CD3803EF2D28CD5C7E3A38E001C00FE2E003EF2D28CD5C7D3A38",
    init_23 => X"2831EF0D4DC324B7CD3803EF2D28CD5C7E3A380103EF2D28CD5C7D3A38010202",
    init_24 => X"310501E5EF2D28CDF5FC3E023004C6FCE606382DD5CD382A0501E50501003234",
    init_25 => X"D5690630B8792307CDC9C13802C31B03A10F31043102C001C11F04A23102C41F",
    init_26 => X"2AC1D9D54F0418C5C1D94F940738BC0338851F78600016D54168C8B107185FAF",
    init_27 => X"4FC50006DF0ACFF328C9D1D91079D922E5CD4F3D0D280D38853C794784785C7D",
    init_28 => X"FE0074CDF32022FE1C8ACA0DFE030074CDE9094E00062684D27916DCCD259621",
    init_29 => X"79190100115C362A2307CDC97E01CBFD1C8AC229FEDF1C79CD062028FEE7C922",
    init_2A => X"1A231407064F3D1A203C0428AE1AE5D5C560065740EE18E6795FA8E0E60F0F0F",
    init_2B => X"2AB2C348D310C1D119000811E10A1812F700010190803EC1C1C1F7100F20A9AE",
    init_2C => X"56A8122BF22E4F281C222D28C37E6758EE03E6796FA8E0E64F0F0F0F792307CD",
    init_2D => X"0FCD1B20250FCD000001E523DF24FFC3E700CEA9C7ABBFAAE6C48FA684A757A5",
    init_2E => X"B6CB5C3B21D10BF22822FE237EF82022FE1312237ED5E1F711282530CDFB2825",
    init_2F => X"764BED28282530CD27BDC32712C3E71C8AC229FE24FBCDE72712C32AB2C47ECB",
    init_30 => X"A77E5C7643ED2DA2CD383103A10232800000418034041637340FA1EF2D2BCD5C",
    init_31 => X"5C3B21270DCA23FEE7105A0126C3C3E73438A3EF04282530CD09187710D60328",
    init_32 => X"010E12F1F7000101F50333CD5F150E30031ECD1320000E028ECD1F287ECBB6CB",
    init_33 => X"CBC42522CD4818E72580C42522CD25DBC3E72535C42522CD2712C32AB2CD0006",
    init_34 => X"230E36231655CD000601DF2C9BCD23202530CD3C3041FE56302C88CD3F18E722",
    init_35 => X"33B4CD23FA200EFE7E23DF0E180077CD2BEBB0ED5C652242EDA7050E5C652AEB",
    init_36 => X"01331833B4CD230438C0FE5C3B3A2996CC1C2EDA28B2CD1418F601CBFD5C5D22",
    init_37 => X"DCC610061C8AD2142814FE04F0011C8ADAAFD62028AEFE10180127282DFE09DB",
    init_38 => X"2A52CD17207601CBFD0C2028FEDF24FFC3E7C5B9CB0238EEFEB1CB0230DFFE4F",
    init_39 => X"3B21C50018CAA73A38B87AD1460926ED214E063016DCCD2795214F0006F018E7",
    init_3A => X"E601AEFD7B0918383BEF473FE67B09282530CDD5991E022076CB0620EDFE7B5C",
    init_3B => X"4F08C63FE615207601CBFD79D5C118C1B6CB02207BCBF6CB5C3B21D11C8AC240",
    init_3C => X"3DC65EC52FC42AC32DCF2B24FFC3E7C5F9CB022817FED7380818F1CB042010FE",
    init_3D => X"2530CD0605050505050503020A08080600C8C6C7C5CBC9CAC8C9C7CD3CCC3ECE",
    init_3E => X"202CFEDF24FBCD102829FEE7122028FEE70120F524FEE71C8AD22C8DCDE73520",
    init_3F => X"204F24D6E747DFE6E72712C3F6CB0228F1B6CB5C3B21E71C8AC229FEF518E703",
    write_mode => "READ_FIRST")
  port map (
    do    => doa(4),
    addr  => addr(10 downto 0),
    clk   => clk,
    en    => ena(4),
    we    => '0',
    ssr   => '0');

  rom5 : RAMB16_S9
  generic map (
    init_00 => X"28ABCD0820B8DFE628ABCDE518CF0230C11D86CDC500CE112B5C532AE5E7E701",
    init_01 => X"FEE528ABCD5C5D53EDD1D128ABCCA7D718C1198BCDC50200112BE10C28B924D6",
    init_02 => X"2B2040E601AEFDF124FBCDD5E52300162328ABCD2B072840160EFE7E23422829",
    init_03 => X"E1E70D202CFEDFE50D2829FE28ABCD2BEBB0ED5C652242ED0005015C652AEBE1",
    init_04 => X"E124FBCDE7E7D55C0B22E35C0B2A5C5D22EBD119CF022829FEDFE5BE1828ABCD",
    init_05 => X"1FE6E51C8AD22C8DCDDFF601CBFDC9FA3821FE7E232712C3E75C0B22E15C5D22",
    init_06 => X"FDE7F618E7B1CB16302C88CD0F302C88CDE9CB112824FEF1CB282828FEE5E74F",
    init_07 => X"5C4B2A37184FFFCBE0E67908202530CD412951C22530CD0628A75C0C3AB601CB",
    init_08 => X"80F6F428BE20F6FA2820FE131A23E5D5D13038293FF287172220B92D287FE67E",
    init_09 => X"D1D10D18E8CB092828FEDFD1F8CBCE18C1EB19B8CDC5E115302C88CD1A0620BE",
    init_0A => X"7E234760F67E28EFCA29FE7E5C0B2AC970CB10CBE1F818E703302C88CDDFE5D1",
    init_0B => X"1828ABCD28EFCA29FE28ABCD23232323231228B978A8CB2328ABCD2B07280EFE",
    init_0C => X"0E207ECB4B2079CB47AFC93CAFD1D15C6522EB33C0CD5C655BED230C2069CBD9",
    init_0D => X"EB612028FEDFEBE828050A2871CB462323232A49C3DF2AB2CDEB2346234E233C",
    init_0E => X"3220CCFE6C2829FEC9E73C2029FE062071CB522879CB20282CFEE1DFE52418EB",
    init_0F => X"2AEECDE5C5E528CCFE512829FEDF0920C0FE79E1E7E50000215E185C5D222BDF",
    init_10 => X"022829FEDF4B42132071CBE5662079CBB310C1D1092AF4CD0B19382ACCCDEBE3",
    init_11 => X"2829FEDF2AB1CDEB4B422309C12AF4CDE32AEECDC9092AF4CD000511E1E702CF",
    init_12 => X"F5AFD5502829FEE72BF1C42530CDC9B601CBFDF82828FEE72A52CDDB202CFE07",
    init_13 => X"186B621C8AC229FE0928CCFEE1DFE55950F52ACDCDF11728CCFEE1DF000111C5",
    init_14 => X"3800000152EDA7E32B19E3F1E62029FE6960DFF52ACDCDF10C2829FEE1E7E513",
    init_15 => X"23775C652AC133A9CDC5B601CBFDAFC82530CDB601CBFDD14D442A20FAA72307",
    init_16 => X"B178D11E99CDF512282530CDF11C82CDF5E5D5AFC95C65222370237123722373",
    init_17 => X"2AC91F15DA30A9CDC82530CDC956235E23EBC9D1E100DE7A42EDA7E5E1052837",
    init_18 => X"CDED18230D3016FE113810FE0B30FA2820FE7E23030005015E284E37CBFD5C4D",
    init_19 => X"7E2311284706D61B5C4D2AD5EB23231655CD2B5C592A792BC0CA24FEE7382C88",
    init_1A => X"0501E13802EFE52BEACDE120F6AE5C4D2AC03E1280F6F410121320F6FA3821FE",
    init_1B => X"7830204637CBFD5C724BED5C4D2AE7181900061106287601CBFD401842EDA700",
    init_1C => X"28B178EBE34D4402300942EDA7E3E12BF1CDE5B8ED2036235D54C5D5F7E5C8B1",
    init_1D => X"19E8C3030303E1C12BC6CDC5E57E2B2B2BC9E1B0EDD5C8B178EBE1D1C1B0ED02",
    init_1E => X"C5C15C4D2A1655CD2B5C592A0303035C4D222BC509EB2BF1CDF5A65C4D2ADF3E",
    init_1F => X"65227E2B5E2B562B4E2B462B5C652AC92B5C592A772BF1712B70C123EBB8ED03",
    init_20 => X"CBC119E8CD19B8CDC508381BEECD2996CDB1CB08202530CD1C8AC228B2CDC95C",
    init_21 => X"2AF4CD6960E524C5E12A20DA2ACCCDFF26E7EB052E022071CB000121C50006F9",
    init_22 => X"2B5C592A4D44E5C5D51F15DA1929232300266879C1E7BB2029FEE8282CFEDFEB",
    init_23 => X"C1B8EDC12036022871CB00361B6B62772378C1702371230B0B0BC177231655CD",
    init_24 => X"111920C4FEC97BFED03F61FED85BFED03F41FED83F2D1BCDC9F8203D2B712B70",
    init_25 => X"FE2D3BCD0F282EFE2D2BC34B42EF18EB31ADDA6AED3FEB0A2000CE31D6E70000",
    init_26 => X"0B382D22CDDF3802C0A1EF38A0EF1C8ADA2D1BCDE70A1822382D1BCDE728202E",
    init_27 => X"CDE70402202DFE05282BFEE7FF06C065FE032845FEEF18E7380F04C005A4E0EF",
    init_28 => X"3AFED830FE2D4FC344ED02280431ADFAA731ADDAC12DD5CD2D3BCDC5CB382D1B",
    init_29 => X"F138A0EFF5C9A738EF2AB6CD4748515FAF5C3A21FD00064F30D6D82D1BCDC93F",
    init_2A => X"F138A4EF350BCD5C9221F53C2F02300F07F1180074CD380F04A401EFD82D22CD",
    init_2B => X"23C93802EFE518F1380431EFF50828F138E1050233040400E0C1EFF50D303FCB",
    init_2C => X"00362377A9897A237791A97B2371230036E5000EC957A9897E235F91A97E234E",
    init_2D => X"E1D17B4B4279CB90AF2D7FCD46EBD5E53802EF38270FA2EF0528A77E38EFC9E1",
    init_2E => X"37F103280405F5D82DA2CD382704859A201AEF34EF2AB6CD47AF4F5F9F1757C9",
    init_2F => X"E5D93802C5C4C3A0EFD72D3E382AC9D7303E38020D0037310B003631EFC9F1C9",
    init_30 => X"D9D50806530928B30620A77A10062D7FCD4720A77E3802C201E203C22731EFD9",
    init_31 => X"38E103C12731EF2D4FCD7A5CAC32925CAC3A572DC1CD7ED67E38E2EF5718D9D1",
    init_32 => X"D62DC1CD13381CFE80D62ECFC3E1778623775CAB213C9F173D5CA132E52DD5CD",
    init_33 => X"D912CB23CB4780D6D97DFACBD92FBACDEB92182D4FCD44ED7877865CAC214707",
    init_34 => X"0E6FED09065CA1115CA621AFE710F8200D2B77278F7E050E5CAA21D912CB13CB",
    init_35 => X"3809D65CAB3AE71023012840CB000E7234FD7134FD13120A200C0D04206FEDFF",
    init_36 => X"FD2FDDCDD9FACB002E95803ED92FBACDEB38E202EF41186FBEFD043E7135FD0A",
    init_37 => X"A121F110C1D9C5572F8BCD7A5F2F8BCD7B0200012018D912CBD9063808FE717E",
    init_38 => X"0528A77700CE7E2BF141090006714EFD5CA121F5D3187134FD7709714EFD795C",
    init_39 => X"09FE785CA1215CAB4BEDD9E1D93802EF7170FD7234FD040136F11008303F0AFE",
    init_3A => X"A779F41015EFCD0D237E0328A7790C18472F52FA90AF15EFCCA72638FCFE0438",
    init_3B => X"3E4F44ED2F83F2A7794AD7453E2F4ACD01061550E61841FB10303ED72E3E04C8",
    init_3C => X"C8A700367EC9D17D4C195929192929545D00266FD51A1BC30006D72B3E02182D",
    init_3D => X"7746234EF5E5C9C179F8107700CE2F7E2B374F4109000501C5C82BFECB7ECB23",
    init_3E => X"FEC8A7C9E1F15E235623D9C1E1D1D9D55E235623D55E57EB46234E23C54E7923",
    init_3F => X"D95D57002EAFD9C03004CDD0C1F2101BCB1ACBD91BCB1ACB2DCBD947C5163021",
    write_mode => "READ_FIRST")
  port map (
    do    => doa(5),
    addr  => addr(10 downto 0),
    clk   => clk,
    en    => ena(5),
    we    => '0',
    ssr   => '0');

  rom6 : RAMB16_S9
  generic map (
    init_00 => X"2356235E23E523D52620B61AEB346ECDEBC9D91401201CD9C014C01CC9000011",
    init_01 => X"93CDD12BC9D12B2B2B72237323779F0B2000CE0F8EEB09EBE146234E237E2323",
    init_02 => X"77E1F12FDDCD2FBACD90F5EB41780330B84F2F9BCDEB472F9BCDE5D5D9E5D932",
    init_03 => X"80E67DD92328342FDDCD013E08301FE1EBD9AD1F6F8D7CEB4AEDEBD9196168E5",
    init_04 => X"CA34D91F073000CE2F7A5F00CE2F7BD95700CE2F7A5F3F44ED7B1F282B7723D9",
    init_05 => X"C9C1F31002381903301711CB0A38290000214D7C1006C53155C3AFD957D931AD",
    init_06 => X"A9CDE14FA9782D7FCD41E3EB2D7FCDD5E5D52220B61AC92BFECBAE23D834E9CD",
    init_07 => X"30C0CDEBD5D9E5D9D830C0CDAF3293CDD1C9D12D8ECD4F0120B37A0A38E1EB30",
    init_08 => X"1DCB1CCBD9D95AEDD919053011182106D962EDE5D962EDA7782FBACDE55A38EB",
    init_09 => X"1F3F173F3DA701208178E1C1D9EBD9EBE4101F19CBD919CB18CBD91DCB1CCBD9",
    init_0A => X"A2D9AF0128803EA77E1530D978D9775C20D97ACBD9063808203CA768303146F2",
    init_0B => X"35D912CB13CBD912CB13CB071220D97ACBD9200629182B77232E3877072FFBCD",
    init_0C => X"1F16CB1778C1D9D5D923E5182834D98016D907203004CD0C3017D718EA10D728",
    init_0D => X"E5D9D830C0CDEBF43830C0CDAFEB3293CD05CFC9D9E1D9D1E173237223712377",
    init_0E => X"D96AEDD929D910CB11CBD911CB171018DF06AF6861D96960E5D92FBACDE5D5D9",
    init_0F => X"28F531D2FA0437D952EDD952EDA70818A7D95AEDD9190F30D952EDD952ED1038",
    init_10 => X"18203E0036063081FEC8A77E313DC39178E1C1D918CBF118CBF15059D9515FE1",
    init_11 => X"303318183E2BFF36237736202BAE803E03202BB62BA6803E2323231A2091FE51",
    init_12 => X"07289000165A043880900806FACB0D01287ACB000E2B2B5E23562391C62FD52C",
    init_13 => X"0036052838CB38CB38CB472BEBD544EDF0A0D67EC9D12D8ECDFA101BCB3ACB47",
    init_14 => X"23AF2D7FCDD5C0A77EEB3296CDC9D1EB77A6FC1027CBFF3E47092807E6FB102B",
    init_15 => X"2B732BEB1DCB1CCB09CBFC302905EB89065853102842B30820A77A9106772B77",
    init_16 => X"CA300F33A1343C368F0A00B040A2DA0F49F100300100B04000B000C9D1702B72",
    init_17 => X"3B353B353B353B352D3014353B353B353B353B353B353B3524351B385131AF30",
    init_18 => X"E23843383337DA37AA37B5367435DE3669346E364534BC35DE359C353B353B35",
    init_19 => X"C6368636A033C0350135C9361F34B334A534AC346A3492384A36AF36C4371337",
    init_1A => X"327835BFCD340F342D341B344932972D4F33A232143783369B34F93506367A33",
    init_1B => X"0E181FE67A6F7CC60F0F0F0F60E6573380F2A7E5237ED95C6553EDD9E3D95C67",
    init_1C => X"664BEDD9D5E333652156235E19002632D7116F07D9095D54FFFB01D9083018FE",
    init_1D => X"C95C6553ED33C0CD5C655BEDC9D1E11F05CD000501E5D5C318D95C673AF1C95C",
    init_1E => X"50C67E2302203FE67E0C4F0707C0E67EC5E3D9E5D933A9CD6B62C9B0ED33A9CD",
    init_1F => X"C8CD000011D5F5C8A7FA181312C805AF47D9E1D9E3C1B0ED0006132391053E12",
    init_20 => X"21E5D96B62C9E133C0CD3406CD5C682AD5C90900064F8107074FF2183DF1D133",
    init_21 => X"4E1A0506C9E1EB33C0CDEB3406CD5C682AEBE5C9D9E1D933C8CD33F7CDD932C5",
    init_22 => X"3362CD33C6CD3803C1E204E031C2A002C00F31335ECD47C9EBF71013237112EB",
    init_23 => X"1F3F17B680E678230B28A77E0006D834E9CD0618FF06C93803E1EE3502C2010F",
    init_24 => X"4F9F2B16CB23000111D5D834E9CDC9D12D8ECD4F2FB178E12D7FCDE5D5C92B77",
    init_25 => X"0B2BF1CDC9C5E52D2B211E99CD2D28C30A1E99CD041878ED1E99CDC9D12D8ECD",
    init_26 => X"815C7B4BED0C30A8FE8787873D3C153015FE193890D609382C8DCD1A2320B178",
    init_27 => X"18FF3ED834E9CDC937C0E1C178B623B623B6237E47C5E509CF2D2BC30401304F",
    init_28 => X"EB34E9CDEBC9E1772377231F771723772377003EE5072BAE23AF051834E9CD06",
    init_29 => X"57CB08D678C9D1121B12AF1BD5D0EB34E9CDEBDE18A7D0EB34E9CDEBE71837D8",
    init_2A => X"C5D52BF1CDF50F3318300FCDF50F072057CBF1EBD1343CCDE5F508300F3D0120",
    init_2B => X"130BED200938961A0D28B11318F116183FF10428C1B10B2078E3B57CE12BF1CD",
    init_2C => X"D52BF1CDC93501D40FF134F9D4F5F13501DCF5F138A0EFF5A7F1C1DF182BE323",
    init_2D => X"2AB0ED0228B178E1C1B0ED0228B178E1C12AB2CDF74D4409C5D5E5E12BF1CDC5",
    init_2E => X"5D2A0ACFC9EB2AB2CD12F1F7000101F50C200E382DD5CDC9D119E5FFFB115C65",
    init_2F => X"24FBCDBE01CBFD0D362BEBB0EDD55C5D53EDE1F703D52BF1CDF59FE3C678E55C",
    init_30 => X"01A0185C5D22E124FBCDFE01CBFD5C5D221C8AC240E601AEFDF1E107200DFEDF",
    init_31 => X"4D4452EDA75C5B2AD11615CDE12DE3CD1601CDFF3EE55C512AE55C5B22F70001",
    init_32 => X"CD12F70C033000000115E6CD1601CDE55C512A1E9FD210FE1E94CDC9EB2AB2CD",
    init_33 => X"355C6721E5D92D2BC32BF1CD2D28C31A0128B1782BF1CD35BFC31615CDE12AB2",
    init_34 => X"C9D9E3D9F1C9D923D9EF20A71B1B1A1313C9D919579F177B5ED9C9D9230420E1",
    init_35 => X"03003001E003C03A31C9383A04003631EFC938E00304C001E02705E03102C0EF",
    init_36 => X"A24065789D66655836138803A10F3103C3273104293BAA38F1343DEFC93803A1",
    init_37 => X"033807202DD5CD38E3CFF87E3AF15894BB7EEE14B0B02FEB24AFF721E7C93260",
    init_38 => X"7E3802A009CF38040037313DEFC938A002EFC97744ED043096073805CF093086",
    init_39 => X"F03401EF34380103A10108003703CDCCCC4CF034310103003834EF2D28CD8036",
    init_3A => X"9EAA905CC53059A5DA560914AC118C03A2042032343103A203A20104F8177231",
    init_3B => X"049380236EF05E7E9CA7ED36CA431BEAFC5CFEA0E7B49F31A496DACBA1616F70",
    init_3C => X"38020400C0373103A12A310F310F3103270FA231046E83F922EE343DEFC9380F",
    init_3D => X"148603A10F3104313139EF03331B0600E003A12A39EFC9381B0200360103A1C9",
    init_3E => X"0520011F31EFC93804EA1B5D23F1EDCD0D92EE23BB6315E9EE388FA30B1F5CE6",
    init_3F => X"0F3104313101A0EF03331B060001A3363105011BA1EF0E3881FE7E3297CDC938",
    write_mode => "READ_FIRST")
  port map (
    do    => doa(6),
    addr  => addr(10 downto 0),
    clk   => clk,
    en    => ena(6),
    we    => '0',
    ssr   => '0');

  rom7 : RAMB16_S9
  generic map (
    init_00 => X"BE3609B5E6C44263B4E8DBA07536009EFD985BBC39588DE4550E13B2108C03A1",
    init_01 => X"3124050FA1281B03A1043131EFC9380F040CB3A161F0BE63DED8EC5D1B7336E9",
    init_02 => X"30310236C4C33804250700303101EF38A21E003031EFC9381B03A322EFC9380F",
    init_03 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC938A1020501A106003701A00900",
    init_04 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_05 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_06 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_07 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_08 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_09 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_0A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_0B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_0C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_0D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_0E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_0F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_10 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_11 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_12 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_13 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_14 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_15 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_16 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_17 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_18 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_19 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_27 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
    init_28 => X"00247E24247E2400000000000024240000100010101010000000000000000000",
    init_29 => X"0000000000100800003A442A102810000046261008646200083E0A3E283E0800",
    init_2A => X"0008083E080800000014083E0814000000201010101020000004080808080400",
    init_2B => X"002010080402000000181800000000000000003E000000001008080000000000",
    init_2C => X"003C42020C423C00007E403C02423C00003E080808281800003C62524A463C00",
    init_2D => X"0010100804027E00003C42427C403C00003C42027C407E0000087E4828180800",
    init_2E => X"20101000001000000010000010000000003C023E42423C00003C42423C423C00",
    init_2F => X"0008000804423C00001008040810000000003E003E0000000004081008040000",
    init_30 => X"003C424040423C00007C42427C427C000042427E42423C00003C405E564A3C00",
    init_31 => X"003C424E40423C00004040407C407E00007E40407C407E000078444242447800",
    init_32 => X"0042444870484400003C424202020200003E080808083E00004242427E424200",
    init_33 => X"003C424242423C000042464A52624200004242425A664200007E404040404000",
    init_34 => X"003C42023C403C000042447C42427C00003C4A5242423C000040407C42427C00",
    init_35 => X"00245A42424242000018244242424200003C424242424200001010101010FE00",
    init_36 => X"000E080808080E00007E201008047E0000101010284482000042241818244200",
    init_37 => X"FF00000000000000001010105438100000701010101070000004081020400000",
    init_38 => X"001C2020201C0000003C22223C202000003C443C04380000007E202078221C00",
    init_39 => X"38043C44443C00000010101018100C00003C407844380000003C44443C040400",
    init_3A => X"0024283030282000182404040400040000381010300010000044444478404000",
    init_3B => X"003844444438000000444444447800000054545454680000000C101010101000",
    init_3C => X"007804384038000000202020201C000006043C44443C00004040784444780000",
    init_3D => X"002854545444000000102828444400000038444444440000000C101010381000",
    init_3E => X"000E080830080E00007C2010087C000038043C44444400000044281028440000",
    init_3F => X"3C4299A1A199423C0000000000281400007010100C1070000008080808080800",
    write_mode => "READ_FIRST")
  port map (
    do    => doa(7),
    addr  => addr(10 downto 0),
    clk   => clk,
    en    => ena(7),
    we    => '0',
    ssr   => '0');
end Behavioral;
