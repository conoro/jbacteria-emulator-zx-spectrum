library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library UNISIM;
use UNISIM.vcomponents.all;

entity vram is port(
    clk     : in  std_logic
  ; rd      : in  std_logic
  ; wr      : in  std_logic
  ; addr    : in  std_logic_vector(13 downto 0)
  ; dataout : out std_logic_vector( 7 downto 0)
);
end vram;

architecture Behavioral of vram is

type EN_a is array(7 downto 0) of std_logic;
type Arr_d is array(7 downto 0) of std_logic_vector(7 downto 0);
signal ENA : EN_a;
signal DOA : Arr_d;

begin

    process(addr, rd, DOA)
    variable i : integer;
    begin
        dataout <= (others => '0');
        for i in 0 to 7 loop
            ENA(i) <= '0';
            if (rd='1' and to_integer(unsigned(addr(13 downto 11))) = i) then
                ENA(i) <= '1';
                dataout <= DOA(i);
            end if;
        end loop;
    end process;

  ram0 : RAMB16_S9
  generic map (
      write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    , INIT_00   => X"9898989898989898989898989898989898989898989898989898989898989898"
    , INIT_01   => X"989800000000000000FF0000FF0000FFFFFFFFFFFF0000000000000000009898"
    , INIT_02   => X"98980003FC01E07FFC01FFC0007FFC00000000000007FFEA8FFF03FFFFE09898"
    , INIT_03   => X"989800FFFFFC000000000000000F000000000000000000000003FFFFF4009898"
    , INIT_04   => X"9898030FFFE0000000000000000000000000000000000000000000FFF9009898"
    , INIT_05   => X"9898003FF0FFFFFFFFFFF800000000000000000000000000000000007F009898"
    , INIT_06   => X"989801FE0001FE00000000000000000000000000001C4768FF80000000309898"
    , INIT_07   => X"989807C000003FC03FF81FFC7E3F1F079F1E7E1E7C3F1F003C3C007E43009898"
    , INIT_08   => X"6262626262626262626262626262626262626262626262626262626262626262"
    , INIT_09   => X"626200000000000000FF0000FF0000FFFFFFFFFFFF8000000000000000006262"
    , INIT_0a   => X"62620007FC03C07FF8007F80007FF000000000000003FF0503FF83FFFFF06262"
    , INIT_0b   => X"626201FFFFF80000000000000006000000000000000000000001FFFFE8006262"
    , INIT_0c   => X"6262070FFFF80000000000000000000000000000000000000000007FFE006262"
    , INIT_0d   => X"6262007FE07FFFFFFFFFF800000000000000000000000000000000001F806262"
    , INIT_0e   => X"626201FC0001FE00000000003780760020003002600E7FFC7FF8000001C06262"
    , INIT_0f   => X"6262078000003FC07FFC1FBC3E3E1E079E1C7F1E7C7F1F00383C00F000C06262"
    , INIT_10   => X"1616161616161616161616161616161616161616161616161616161616161616"
    , INIT_11   => X"161600000000000000FF0000FF0000FFFFFFFFFFFF8000000000000000001616"
    , INIT_12   => X"1616000FFE07C03FE0001F00007FE000000000000000FC0001FFC7FFFFF81616"
    , INIT_13   => X"161601FFFFF80000000000000002000000000000000000000000FFFFD0001616"
    , INIT_14   => X"1616040FFFFE01C0000F40000000000000000000000000000000003FFD001616"
    , INIT_15   => X"1616007FE01FFFFFFFFFF000000000000000000000000000000000000F801616"
    , INIT_16   => X"161601FC0001FF00070033D83FD07FE1383E7003380E7FFE7FF800000F001616"
    , INIT_17   => X"1616078000003FC0FFFC3E1E3E1F1E079E1C3F9E3E3E3F00187C018000301616"
    , INIT_18   => X"BCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBC"
    , INIT_19   => X"BCBC000000000C0000FF0000FF0001FF0FFFFFFFFF000000000000000000BCBC"
    , INIT_1a   => X"BCBC001FFF0F803FC0000400007FC000000000000000300000FFE7FFFFFCBCBC"
    , INIT_1b   => X"BCBC01FFFFF000000000000000000000000000000000000000003FFFE800BCBC"
    , INIT_1c   => X"BCBC001FFEFF8BF8F5DFE0000000000000000000000000000000001FFC80BCBC"
    , INIT_1d   => X"BCBC007FC007FFEFFF81F000000000000000000000000000000000000780BCBC"
    , INIT_1e   => X"BCBC03F80000FF001F807FF87FF83FFFBE3CF80F3C1C3FFC7FFC00007F00BCBC"
    , INIT_1f   => X"BCBC070000003FC0FFFC3C1E3E1F3F070E1E7F9C1FBC3FC01C7C00000008BCBC"
    , INIT_20   => X"A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3"
    , INIT_21   => X"A3A3000000001A0000FF0001FFC000FC00FFFFFFC3000000000000000000A3A3"
    , INIT_22   => X"A3A3003FFF9F001F80000000007FC0000000000000000000007FFFFFFFE4A3A3"
    , INIT_23   => X"A3A301EFFFE000000000000000000000000000000000000000001FFFF400A3A3"
    , INIT_24   => X"A3A3001FFDFFFFFFFFFFE00000000000000000000000000000000007FF00A3A3"
    , INIT_25   => X"A3A300FF8001FF00D60180000000000000000000000000000000000003C0A3A3"
    , INIT_26   => X"A3A303F000007F000FC03FF87FFC3FFF0E3CF80F3C1E3FFE3FFE0001FF00A3A3"
    , INIT_27   => X"A3A30A0000007FC07F7E7C1C1E1C3E071E3E7F1E1F8C3FC03CF800000038A3A3"
    , INIT_28   => X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D"
    , INIT_29   => X"0D0D000000003C0000BF0006C14000F00007FFF002C00000000001FFFE000D0D"
    , INIT_2a   => X"0D0D007FFFBF000F00000000003F80000000000000000000003FFFFFFF280D0D"
    , INIT_2b   => X"0D0D03CFFFE000000000000000000000000000000000000000000FFFF8000D0D"
    , INIT_2c   => X"0D0D001FFFFFFFFFFFFFF80000000000000000000000000000000003FE800D0D"
    , INIT_2d   => X"0D0D00FF8000FE00000000000000000000000000000000000000000001C00D0D"
    , INIT_2e   => X"0D0D03F000007F801FE03FF87FFE3FFF0E3C7C1F1C1E3FFE3EFC0007FF000D0D"
    , INIT_2f   => X"0D0D0A000000FFC0FC3E7C0C1E1C3E1E1E3C7F9E3FCE1FE07DF0000000700D0D"
    , INIT_30   => X"6161616161616161616161616161616161616161616161616161616161616161"
    , INIT_31   => X"6161000000007A00010F0008424000C000007C00012000067FFC01FFFF006161"
    , INIT_32   => X"616100FFFFFE000E00000000001F80000000000000000000000FFFFFFD506161"
    , INIT_33   => X"6161038FFFC0000000000000000000000000000000000000000007FFF4006161"
    , INIT_34   => X"6161003FFDFFFFFFFFFFF80000000000000000000000000000000001FF006161"
    , INIT_35   => X"616100FF00007E00000000000000000000000000000000000000000000406161"
    , INIT_36   => X"616103E000007F803FF01FFE3FFF3FFF1C3E7E0E1C1E1FFA1C7E000FFF006161"
    , INIT_37   => X"61610C000000FF80F81E1E0C1E3E7E3C1C3EFFDF3FCF1FF07FF0000000F06161"
    , INIT_38   => X"3232323232323232323232323232323232323232323232323232323232323232"
    , INIT_39   => X"323200007800F400020300320040030000000000001800181FFE03FFFF003232"
    , INIT_3a   => X"323200FFFFFE000400000000000F000000000000000000000007FFFFFA803232"
    , INIT_3b   => X"3232038FFFC0000000000000000000000000000000000000000003FFFA003232"
    , INIT_3c   => X"3232003FFAFFFFFFFFFFF00000000000000000000000000000000000FF003232"
    , INIT_3d   => X"323201FF0000FE0000000000000000000000000000000000E180000000203232"
    , INIT_3e   => X"323207E000003F803FF81FFC7FFE1E3F0F1E3E1C3C1E1F801C3E001FCF003232"
    , INIT_3f   => X"32320C000001FF01F81F1E1C1E3E7E7C1E0E3FDF3FFF1FF03F80000003E03232"
  )
  port map (
      DI    => "00000000"
    , DIP   => "0"
    , DO    => DOA(0)
    , ADDR  => addr(10 downto 0)
    , CLK   => clk
    , EN    => ENA(0)
    , WE    => '0'
    , SSR   => '0'
  );

  ram1 : RAMB16_S9
  generic map (
      write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    , INIT_00   => X"9898F8000001FF01F03E1E1E3F3E7FF00E0E3FFE1FFE1FF07F80000007E09898"
    , INIT_01   => X"9898F0000000FF803FF07E1F07FC3EFE1FFE383F7F0F3FDC1E1F003FFF009898"
    , INIT_02   => X"9898E00000000000000000000000000000000000000000000001FFFFE0009898"
    , INIT_03   => X"9898FF000080C000000000000000000000000000000000000FFFFFFC00009898"
    , INIT_04   => X"9898F00001023CFFBC00000200000000000000000000007FFFFFFF8000009898"
    , INIT_05   => X"9898F8000053FFFFFF00000F08042110000000000007FFFFFFFFF80000009898"
    , INIT_06   => X"989850001A871FFE00EA000000000000010000003FFFFFFFEFFFF80000009898"
    , INIT_07   => X"98983EA000F0BF410040F00000000000000001FFF0000000003FF00000009898"
    , INIT_08   => X"6262F0000001FE00F87E1F3F3F3C3FF00E1E73FE3DFF1FC07FF000001FE06262"
    , INIT_09   => X"6262F80000007F801FF83E1F87F83E3F0FFC383E7F0F1FFC1E1F00FFFE006262"
    , INIT_0a   => X"6262F00000006000000000000000000000000000000000000007FFFFC0006262"
    , INIT_0b   => X"6262FE000080D800000000000000000000000000000000003FFFFFF800006262"
    , INIT_0c   => X"6262F8000104427F42C000020003008400000000000001FFFFFFFF8000006262"
    , INIT_0d   => X"6262F00000A3FEF7FF008000100421138EE31C00000FFFFFFFFFF80000006262"
    , INIT_0e   => X"62626800148300000050000000000000010000007FFFC0FFC7FFF80000006262"
    , INIT_0f   => X"62623F5000F8BF000020F00000000000000003FFF0000000007FF00000006262"
    , INIT_10   => X"1616F0000001FE00FCFE1FFF0F3E3FF00E3E73FE3CFF3E003FF000003FC01616"
    , INIT_11   => X"1616F80000007F000FF03E0F0FF03E7E0FFC781E7F0F0FFC1E1E01FFFE001616"
    , INIT_12   => X"1616FC000001C00000000000000000000000000000000000000FFFFFC0001616"
    , INIT_13   => X"1616F8000000F800000000000000000000000000000000007FFFFFF800001616"
    , INIT_14   => X"1616F8000005F11C8FE000040002C08800000000000003FFFFFFFF0000001616"
    , INIT_15   => X"1616F00000A7FFFFFF008000200442249094A000001FFFFFFFFFF80000001616"
    , INIT_16   => X"161674002F800000018E00000000000001000000FFFF807F07FFF80000001616"
    , INIT_17   => X"16163FB000F8BF000020F8000000000000000FFFE000000000FFF00000001616"
    , INIT_18   => X"BCBCE0000001FE01FFFF1FFF3F3E3FF80C3E70FE1C7E3E003FF000007FC0BCBC"
    , INIT_19   => X"BCBCFC0000007E0007F03C0F8FF07E0F1FFCF80F3E031FFF8C0703FFFC00BCBC"
    , INIT_1a   => X"BCBCFE000007C00000000000000000000000000000000000001FFFFF8000BCBC"
    , INIT_1b   => X"BCBCF0000000A80000000000000000000000000000000001FFFFFFF00000BCBC"
    , INIT_1c   => X"BCBCF800000ABD42BD500004000220880000000000000FFFFFFFFF000000BCBC"
    , INIT_1d   => X"BCBCE000014783F87F00C0004004422490972000007FFFFFFFFFF8000000BCBC"
    , INIT_1e   => X"BCBC3A002F80F0000F3F00000000000002000003FFFF807E03FFF8000000BCBC"
    , INIT_1f   => X"BCBC1FD8007DBF000050F8000000000000001FFFE000000001FFE0000000BCBC"
    , INIT_20   => X"A3A3C0000001FE00FFFE1FFF9F3E3FF80E3E307F1C7E1E007FFE0001FF80A3A3"
    , INIT_21   => X"A3A3FC0000007E0003C0380F8FF0740F1FFCF80F3C03BF871C030FFFFC00A3A3"
    , INIT_22   => X"A3A3FF00000FC00000000000000000000000000000000000007FFFFF8000A3A3"
    , INIT_23   => X"A3A3E0000000AC0000000000000000000000000000000003FFFFFFE00000A3A3"
    , INIT_24   => X"A3A3FC000016FF24FE580004000220880000000000001FFFFFFFFE000000A3A3"
    , INIT_25   => X"A3A3E000078200E01F0CC010800482249094200000FFFFFFFFFFF8000000A3A3"
    , INIT_26   => X"A3A33D0053C0CFFFF0FF80000000000000000007FDFF003C01FFF8000000A3A3"
    , INIT_27   => X"A3A31FF4007FBF000028FC000000000000003FFFC000000003FFE0000000A3A3"
    , INIT_28   => X"0D0DE0000001FE007FFC1FFF0F3E1FFF0E3C703F3C7F1F003FFE0003FF800D0D"
    , INIT_29   => X"0D0DF80000003C0000007800000000001000200230039F001C001FFFF8000D0D"
    , INIT_2a   => X"0D0DFF80001F80000000000000000000000000000000000000FFFFFF00000D0D"
    , INIT_2b   => X"0D0DE00001005F0000000000000000000000000000000007FFFFFFE000000D0D"
    , INIT_2c   => X"0D0DFC00001239009C5C000B220210880000000000003FFFFFFFFE0000000D0D"
    , INIT_2d   => X"0D0DC0000EC00000077080130007122350E3A10001FFFFFFFFFFF80000000D0D"
    , INIT_2e   => X"0D0D3A0063C0800000FFC000000000000000001FFC00001000FFF80000000D0D"
    , INIT_2f   => X"0D0D1FFA003FBF000018FC00000000000000FFFFC0000001C7FFE00000000D0D"
    , INIT_30   => X"6161E0000001FF003FF83F3F0FFC3EFF1F7C783F3E1F1F007E7E0007FF806161"
    , INIT_31   => X"6161E00000003C000000000000000000000000000000000000007FFFF0006161"
    , INIT_32   => X"6161FFC0003F80000000000000000000000000000000000003FFFFFE00006161"
    , INIT_33   => X"6161F000011841000000000000000000000000000000001FFFFFFFC000006161"
    , INIT_34   => X"6161FC00002B860061E6000892021110000000000000FFFFFFFFFC0000006161"
    , INIT_35   => X"6161E0000F8000000081800C000000000080000007FFFFFFFFFFF80000006161"
    , INIT_36   => X"61613D8001E0810040FFC000000000000000003FF800000000FFF00000006161"
    , INIT_37   => X"61611FF5003FDF000024FE00000000000001FFFFC0000000BFFF800000006161"
    , INIT_38   => X"3232F0000000FF003FF87E1F0FFC1E7E1FFE783F7F0E1F001E3F001FFF003232"
    , INIT_39   => X"3232C00000001800000000000000000000000000000000000000FFFFF0003232"
    , INIT_3a   => X"3232FF80003F80000000000000000000000000000000000007FFFFFE00003232"
    , INIT_3b   => X"3232F000017E7E003C00000200000000000000000000003FFFFFFFC000003232"
    , INIT_3c   => X"3232F80000517C003EFF0008940411F0000000000001FFFFFFFFFC0000003232"
    , INIT_3d   => X"3232E0001F0400000702000000000000010000000FFFFFFFFFFFF80000003232"
    , INIT_3e   => X"32323F4001E0208080FFE000000000000000007FF8000000007FF00000003232"
    , INIT_3f   => X"32320FFB001F9F000016FF00000000000003FFFFC00000007FFC000000003232"
  )
  port map (
      DI    => "00000000"
    , DIP   => "0"
    , DO    => DOA(1)
    , ADDR  => addr(10 downto 0)
    , CLK   => clk
    , EN    => ENA(1)
    , WE    => '0'
    , SSR   => '0'
  );

  ram2 : RAMB16_S9
  generic map (
      write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    , INIT_00   => X"989807FD800F0F42000B008000000000000FFFFFC00000003FF0000000009898"
    , INIT_01   => X"9898007FF50000E00000AFFF00000000FFFC0000000000000000000000009898"
    , INIT_02   => X"989801FFFFF4000000000100700003FFFFE00000000000000000000000009898"
    , INIT_03   => X"9898007FC00750370702555F081FFFF800000000000000000000003FFC009898"
    , INIT_04   => X"98980018007FFEA003C003FFFFE0FFFFE0007FFDDF77FFFFF7DCFFFFFFFF9898"
    , INIT_05   => X"98980000001F00FEAD45AFE00000000000007EC1DB77E49554503FFC3FFC9898"
    , INIT_06   => X"9898989898989898989898989898989898989898989898989898989898989898"
    , INIT_07   => X"9898989898989898989898989898989898989898989898989898989898989898"
    , INIT_08   => X"626201FF40060081F80780C000000000001FFFFFC00000001F80000000006262"
    , INIT_09   => X"6262007FFB0000F03F001F7F00000001FFF80000000000000000000000006262"
    , INIT_0a   => X"626201FFFFFA000C00000100780007FFFFC00000000000000000000000006262"
    , INIT_0b   => X"6262007E8007E80A0301A0AF043FFFF800000000007000000F70000FE0006262"
    , INIT_0c   => X"62620018007FFF6001E000FFFFC0FFFFF80000000070000014503FFC3FFC6262"
    , INIT_0d   => X"62620000001E003F7D875FC00000000000006EC1DB76E255545007E007E06262"
    , INIT_0e   => X"6262626262626262626262626262626262626262626262626262626262626262"
    , INIT_0f   => X"6262626262626262626262626262626262626262626262626262626262626262"
    , INIT_10   => X"161600FFA0000700000BC0C000000000007FFF9FC00000000C00000000001616"
    , INIT_11   => X"1616007FFD8000FFC0E0073F80000003FFFC2493ABB0A9A8CECE4C8924CE1616"
    , INIT_12   => X"161601FFFFF40003200001007C001FFFFF806623624476244000000000001616"
    , INIT_13   => X"1616007F000FF4038100505700FFFFF800000000007000001150000180001616"
    , INIT_14   => X"16160010003FFFB000F8003EFF807FFFFE00000000700000145007E007E01616"
    , INIT_15   => X"161600000018000FAA04BF000000000000006EC1DB76E1555450018001801616"
    , INIT_16   => X"1616161616161616161616161616161616161616161616161616161616161616"
    , INIT_17   => X"1616161616161616161616161616161616161616161616161616161616161616"
    , INIT_18   => X"BCBC007F500003000005F0E00000000000FFFF01C0000000000000000000BCBC"
    , INIT_19   => X"BCBC007FFF4000F00018031FC0000007FFF854A92A28AA28A8A8AADAA528BCBC"
    , INIT_1a   => X"BCBC01FFFFFB8000D400020036003EFBFF005554556C4556C00000000000BCBC"
    , INIT_1b   => X"BCBC007F001FEA004100A80B01FFFFF80000000000700000175000000000BCBC"
    , INIT_1c   => X"BCBC0000003FFFE8007C001D80003FFFFF003CB9CE73C7C7145001800180BCBC"
    , INIT_1d   => X"BCBC000000100003F4035C000000000000006EC1DF76EF52545C00000000BCBC"
    , INIT_1e   => X"BCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBC"
    , INIT_1f   => X"BCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCAC"
    , INIT_20   => X"A3A3001FB00001110002F8F00000000001FFFC0000000000000000000000A3A3"
    , INIT_21   => X"A3A300FFFFA000000004030FC000000FFFFC56A92A28AA28A8A8AAAAB508A3A3"
    , INIT_22   => X"A3A300FFFEF5C0002A8003802B00FFF8FE00555455544555400000018000A3A3"
    , INIT_23   => X"A3A3003E001FF600A000D00707FFFFF80000000000700000145000000000A3A3"
    , INIT_24   => X"A3A30000003FFFF4002B002E0000000000007EFDDF77E848945000000000A3A3"
    , INIT_25   => X"A3A30000000000003803E8000000000000007EC1DF77E848944400000000A3A3"
    , INIT_26   => X"A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3"
    , INIT_27   => X"A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3FF"
    , INIT_28   => X"0D0D001FD800001080017CF80000000007FFF800000000000000000000000D0D"
    , INIT_29   => X"0D0D00FFFF501F0000000107E000003FFFF875A93B30EAB8CCCCAC8BAD0C0D0D"
    , INIT_2a   => X"0D0D00FFFC3A7500155006403581FFF87E0066556744665440000007E0000D0D"
    , INIT_2b   => X"0D0D003E003FFB00C000E8010FFFFFF800007FFDDF77FFFFF7DC018001800D0D"
    , INIT_2c   => X"0D0D0000003FFFEA0035801500000000000066CDDF766BD25450000000000D0D"
    , INIT_2d   => X"0D0D0000000000000803800000000000000036C1CE736F871C7C000000000D0D"
    , INIT_2e   => X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D"
    , INIT_2f   => X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0EE0"
    , INIT_30   => X"6161003FF40000A04002BEFC000000000FFFF000000000000000000000006161"
    , INIT_31   => X"616100FFFFB07F0000000101E000007FFFF054A92A28AAA888A8AA8AA5286161"
    , INIT_32   => X"616100FFF80DBC800FA81D803683FFF83C004555554445544CCC003FFC006161"
    , INIT_33   => X"6161003C003FFE80E080F0001FFBFFFE00004005D1740000000407E007E06161"
    , INIT_34   => X"61610000003FEFF6001AC02A0000000000000EC1DB70EA155450000000006161"
    , INIT_35   => X"6161000000000000000000000000000000000000000000000000000000006161"
    , INIT_36   => X"6161616161616161616161616161616161616161616161616161616161616161"
    , INIT_37   => X"61616161616161616161616161616161616161616161616161616161616162EA"
    , INIT_38   => X"3232003FFA0000C000015EFE000000003FFF0000000000000000000000003232"
    , INIT_39   => X"323200FFFFD8FF0000000100F00001FFFFE054912BA8A9A88EA84A8AA4CE3232"
    , INIT_3a   => X"323200FFE0025F5007FFEA601B0FFFF808004523554445244CCC00FFFF003232"
    , INIT_3b   => X"3232003C007FFD40F880F8007FF1FFFF80004005D174000000043FFC3FFC3232"
    , INIT_3c   => X"32320000003F837B082B01550000000000003EC1DB73E9155450000000003232"
    , INIT_3d   => X"3232000000000000000000000000000000000000000000000000000000003232"
    , INIT_3e   => X"3232323232323232323232323232323232323232323232323232323232323232"
    , INIT_3f   => X"323232323232323232323232323232323232323232323232323232323232322A"
  )
  port map (
      DI    => "00000000"
    , DIP   => "0"
    , DO    => DOA(2)
    , ADDR  => addr(10 downto 0)
    , CLK   => clk
    , EN    => ENA(2)
    , WE    => '0'
    , SSR   => '0'
  );

  ram3 : RAMB16_S9
  generic map (
      write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    , INIT_00   => X"7878787878787878787878787878787878787878787878787878787878787878"
    , INIT_01   => X"78780A0A0A0A0A0A09010A09010909010101010101090A090A0A0A0A0A0A7878"
    , INIT_02   => X"78780A0A0A0A02010101010102010102020202020201010101020A0A0A0A3878"
    , INIT_03   => X"78780A0A0A020202020202020201020202020202020202020202020A0A0A3878"
    , INIT_04   => X"78780A0A3246464646464602020202020202020202020202020202020A0A3878"
    , INIT_05   => X"78780A0A024646464646460202020202020202020202020206060202020A3878"
    , INIT_06   => X"78780A0202064606464646464646464646464646464646464646020101093878"
    , INIT_07   => X"78780A0202064646464646464646464646464646464646464646010101093878"
    , INIT_08   => X"78780102024646064646464646464646464646464646464646460602020A3878"
    , INIT_09   => X"7878010202024646464646464646464646464646464646464646020A0A0A3878"
    , INIT_0a   => X"78780101434343030202024242424242424202020202020202020A0A0A0A3878"
    , INIT_0b   => X"787801020358430304030242424242424242020202020202020A0A0A0A0A3878"
    , INIT_0c   => X"78780102430484202004034242454545424202020202020A0A0A0A0A0A0A3878"
    , INIT_0d   => X"7878010204040C0C0C200442424545454545450202020A0A0A0A0A0A0A0A3878"
    , INIT_0e   => X"78780A02040420202004044242424242454202020A0A0A0A0A0A0A0A0A0A3878"
    , INIT_0f   => X"78780A020304042020200402020202020202020A0A0A0A0A0A0A0A0A0A0A3878"
    , INIT_10   => X"78780A0A02440420202020040202020202020A0A0A0A0A0A0A0A0A0A0A0A3878"
    , INIT_11   => X"78780A0A0202042020202004040202020A0A4747474747474747474747473878"
    , INIT_12   => X"78780A0A0A0A2020202020040402020A0A0A4747474747474747464141463878"
    , INIT_13   => X"78780A0A0A0A02042004202002020A0A0A0A4747474747474747415121413878"
    , INIT_14   => X"78780A0A0A0A0A02040404040A0A0A0A0A0A4747474747474747512151213878"
    , INIT_15   => X"78780A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A4747474747474747420442043878"
    , INIT_16   => X"7878783838383838383838383838383838383838383838383838383838383878"
    , INIT_17   => X"7878787878787878787878787878787878787878787878787878787878787878"
  )
  port map (
      DI    => "00000000"
    , DIP   => "0"
    , DO    => DOA(3)
    , ADDR  => addr(10 downto 0)
    , CLK   => clk
    , EN    => ENA(3)
    , WE    => '0'
    , SSR   => '0'
  );

    RAMB : for i in 4 to 7 generate
    RAMB16_S9_inst : RAMB16_S9
    generic map (
        write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    )
    port map (
        DO => DOA(i),      -- 8-bit Data Output
        ADDR => addr(10 downto 0),  -- 11-bit Address Input
        CLK => clk,    -- Clock
        DI => "00000000",      -- 8-bit Data Input
        DIP => "0",
	     EN => ENA(i),      -- RAM Enable Input
        SSR => '0',    -- Synchronous Set/Reset Input
        WE => '0'       -- Write Enable Input
    );
    end generate;

--  ram4 : RAMB16_S9
--  generic map (
--      write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
--  )
--  port map (
--      DI    => "00000000"
--    , DO    => dataout
--    , ADDR  => "00000000000"
--    , CLK   => clk
--    , EN    => ram4en
--    , WE    => '0'
--    , SSR   => '0'
--  );

end Behavioral;
