library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ram is port(
    clk   : in  std_logic;
    wr    : in  std_logic;
    addr  : in  std_logic_vector(13 downto 0);
    din   : in  std_logic_vector( 7 downto 0);
    dout  : out std_logic_vector( 7 downto 0));
end ram;

architecture behavioral of ram is

  type ram_t is array (0 to 16383) of std_logic_vector(7 downto 0);
  signal ram : ram_t := (
  X"E7", X"DF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --0000
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --0008
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FC", X"00", --0010
  X"00", X"00", X"00", X"00", X"00", X"00", X"3F", X"FF", --0018
  X"FF", X"DF", X"FF", X"FF", X"80", X"7F", X"F0", X"00", --0020
  X"00", X"01", X"8F", X"FF", X"FF", X"FF", X"FF", X"FF", --0028
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"81", --0030
  X"01", X"00", X"00", X"00", X"00", X"80", X"FF", X"FF", --0038
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0040
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0048
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0050
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0058
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0060
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0068
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0070
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0078
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0080
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0088
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0090
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0098
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --00A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --00A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --00B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --00B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --00C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --00C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --00D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --00D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --00E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --00E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --00F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --00F8
  X"81", X"BF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --0100
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --0108
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F8", X"00", --0110
  X"00", X"00", X"00", X"00", X"00", X"00", X"0F", X"FF", --0118
  X"6D", X"EF", X"FF", X"FC", X"00", X"07", X"E0", X"00", --0120
  X"00", X"00", X"73", X"FF", X"FF", X"FF", X"FF", X"FF", --0128
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"E3", --0130
  X"03", X"80", X"1C", X"0E", X"03", X"C1", X"FF", X"FF", --0138
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0140
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0148
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0150
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0158
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0160
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0168
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0170
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0178
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0180
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0188
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0190
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0198
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --01A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --01A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --01B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --01B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --01C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --01C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --01D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --01D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --01E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --01E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --01F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --01F8
  X"01", X"F9", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --0200
  X"FF", X"F1", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --0208
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F8", X"00", --0210
  X"00", X"00", X"00", X"00", X"00", X"00", X"03", X"FF", --0218
  X"EE", X"FF", X"FF", X"F0", X"00", X"00", X"F0", X"00", --0220
  X"00", X"00", X"0F", X"7F", X"FF", X"FF", X"FF", X"FF", --0228
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --0230
  X"87", X"80", X"3E", X"1F", X"8F", X"E3", X"FF", X"FF", --0238
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0240
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0248
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0250
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0258
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0260
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0268
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0270
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0278
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0280
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0288
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0290
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0298
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --02A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --02A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --02B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --02B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --02C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --02C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --02D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --02D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --02E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --02E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --02F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --02F8
  X"00", X"C7", X"FF", X"FF", X"FF", X"FF", X"FF", X"FC", --0300
  X"3F", X"C0", X"7F", X"FF", X"FF", X"FF", X"FF", X"FF", --0308
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F8", X"00", --0310
  X"00", X"00", X"00", X"00", X"00", X"00", X"03", X"FF", --0318
  X"DE", X"FF", X"FF", X"E0", X"00", X"00", X"0F", X"E0", --0320
  X"00", X"00", X"00", X"7F", X"FF", X"FF", X"E0", X"00", --0328
  X"03", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --0330
  X"FF", X"F8", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --0338
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0340
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0348
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0350
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0358
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0360
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0368
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0370
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0378
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0380
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0388
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0390
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0398
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --03A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --03A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --03B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --03B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --03C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --03C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --03D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --03D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --03E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --03E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --03F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --03F8
  X"00", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"C0", --0400
  X"03", X"C0", X"7F", X"FF", X"FF", X"FF", X"FF", X"FF", --0408
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FC", X"00", --0410
  X"00", X"00", X"00", X"00", X"00", X"00", X"03", X"FF", --0418
  X"DE", X"FF", X"FF", X"C0", X"00", X"00", X"00", X"1F", --0420
  X"F0", X"00", X"00", X"01", X"FF", X"F0", X"00", X"00", --0428
  X"00", X"07", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --0430
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F0", --0438
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0440
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0448
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0450
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0458
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0460
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0468
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0470
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0478
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0480
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0488
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0490
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0498
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --04A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --04A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --04B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --04B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --04C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --04C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --04D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --04D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --04E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --04E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --04F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --04F8
  X"80", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", --0500
  X"00", X"30", X"3F", X"FF", X"FF", X"FF", X"FF", X"FF", --0508
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"80", --0510
  X"00", X"00", X"00", X"00", X"00", X"00", X"03", X"FF", --0518
  X"DF", X"7F", X"FF", X"80", X"00", X"00", X"00", X"00", --0520
  X"00", X"00", X"00", X"00", X"00", X"0F", X"E0", X"00", --0528
  X"00", X"00", X"1F", X"FF", X"FF", X"FF", X"FF", X"FF", --0530
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"C0", --0538
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0540
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0548
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0550
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0558
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0560
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0568
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0570
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0578
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0580
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0588
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0590
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0598
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --05A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --05A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --05B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --05B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --05C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --05C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --05D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --05D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --05E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --05E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --05F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --05F8
  X"80", X"FF", X"FF", X"FF", X"FF", X"FF", X"FE", X"00", --0600
  X"00", X"0C", X"3F", X"FF", X"FF", X"FF", X"FF", X"FF", --0608
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"80", --0610
  X"00", X"00", X"00", X"00", X"00", X"00", X"07", X"FF", --0618
  X"FF", X"FF", X"FE", X"00", X"00", X"00", X"00", X"00", --0620
  X"00", X"00", X"00", X"00", X"00", X"00", X"0F", X"FF", --0628
  X"00", X"00", X"00", X"00", X"3F", X"FF", X"FF", X"FF", --0630
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"80", --0638
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0640
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0648
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0650
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0658
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0660
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0668
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0670
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0678
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0680
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0688
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0690
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0698
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --06A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --06A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --06B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --06B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --06C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --06C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --06D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --06D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --06E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --06E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --06F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --06F8
  X"C3", X"BF", X"FF", X"FF", X"FF", X"FF", X"F8", X"00", --0700
  X"00", X"02", X"1F", X"FF", X"FF", X"FF", X"FF", X"FF", --0708
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"80", --0710
  X"00", X"00", X"00", X"00", X"00", X"00", X"0F", X"FF", --0718
  X"FF", X"FF", X"F8", X"00", X"00", X"00", X"00", X"00", --0720
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0728
  X"00", X"00", X"00", X"00", X"00", X"03", X"FF", X"FF", --0730
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", --0738
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0740
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0748
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0750
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0758
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0760
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0768
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0770
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0778
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0780
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0788
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0790
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0798
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --07A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --07A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --07B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --07B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --07C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --07C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --07D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --07D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --07E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --07E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --07F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --07F8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0800
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0808
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"3C", --0810
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0818
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0820
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0828
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0830
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0838
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0840
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0848
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0850
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0858
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0860
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0868
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0870
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0878
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0880
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0888
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0890
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0898
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --08A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --08A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --08B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --08B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --08C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --08C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --08D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --08D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --08E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --08E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --08F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --08F8
  X"00", X"42", X"00", X"42", X"7C", X"00", X"00", X"00", --0900
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0908
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"42", --0910
  X"00", X"7C", X"42", X"40", X"40", X"3C", X"7C", X"00", --0918
  X"00", X"42", X"00", X"78", X"3C", X"42", X"42", X"00", --0920
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0928
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0930
  X"00", X"00", X"18", X"3C", X"3C", X"08", X"00", X"00", --0938
  X"00", X"7E", X"00", X"40", X"7E", X"7E", X"FE", X"00", --0940
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0948
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0950
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0958
  X"00", X"42", X"00", X"7C", X"3E", X"3C", X"42", X"FE", --0960
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0968
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0970
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0978
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0980
  X"00", X"00", X"00", X"3C", X"3C", X"3C", X"7C", X"7E", --0988
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0990
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0998
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --09A0
  X"00", X"00", X"00", X"42", X"3E", X"3C", X"42", X"00", --09A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --09B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --09B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --09C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --09C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --09D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --09D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --09E0
  X"00", X"00", X"3C", X"7C", X"3C", X"3C", X"7E", X"00", --09E8
  X"FE", X"3C", X"00", X"3C", X"FE", X"3C", X"7C", X"FE", --09F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --09F8
  X"00", X"62", X"00", X"42", X"42", X"00", X"00", X"00", --0A00
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0A08
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"99", --0A10
  X"00", X"42", X"42", X"40", X"40", X"42", X"42", X"00", --0A18
  X"00", X"66", X"00", X"44", X"42", X"42", X"62", X"00", --0A20
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0A28
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0A30
  X"00", X"00", X"28", X"42", X"42", X"18", X"00", X"00", --0A38
  X"00", X"04", X"00", X"40", X"40", X"40", X"10", X"00", --0A40
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0A48
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0A50
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0A58
  X"00", X"24", X"00", X"42", X"08", X"42", X"42", X"10", --0A60
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0A68
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0A70
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0A78
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0A80
  X"00", X"00", X"00", X"40", X"42", X"42", X"42", X"40", --0A88
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0A90
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0A98
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0AA0
  X"00", X"00", X"00", X"42", X"08", X"42", X"42", X"00", --0AA8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0AB0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0AB8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0AC0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0AC8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0AD0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0AD8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0AE0
  X"00", X"00", X"40", X"42", X"42", X"42", X"40", X"00", --0AE8
  X"10", X"42", X"00", X"40", X"10", X"42", X"42", X"10", --0AF0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0AF8
  X"00", X"52", X"00", X"42", X"42", X"00", X"00", X"00", --0B00
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0B08
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"A1", --0B10
  X"00", X"7C", X"42", X"40", X"40", X"42", X"42", X"00", --0B18
  X"00", X"5A", X"00", X"42", X"42", X"42", X"52", X"00", --0B20
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0B28
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0B30
  X"00", X"00", X"08", X"42", X"3C", X"28", X"00", X"00", --0B38
  X"00", X"08", X"00", X"40", X"7C", X"7C", X"10", X"00", --0B40
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0B48
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0B50
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0B58
  X"00", X"18", X"00", X"42", X"08", X"40", X"7E", X"10", --0B60
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0B68
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0B70
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0B78
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0B80
  X"00", X"00", X"00", X"3C", X"40", X"42", X"42", X"7C", --0B88
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0B90
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0B98
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0BA0
  X"00", X"00", X"00", X"7E", X"08", X"40", X"7E", X"00", --0BA8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0BB0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0BB8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0BC0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0BC8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0BD0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0BD8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0BE0
  X"00", X"00", X"3C", X"42", X"42", X"40", X"7C", X"00", --0BE8
  X"10", X"42", X"00", X"3C", X"10", X"42", X"42", X"10", --0BF0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0BF8
  X"00", X"4A", X"00", X"42", X"7C", X"00", X"00", X"00", --0C00
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0C08
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"A1", --0C10
  X"00", X"42", X"42", X"40", X"40", X"7E", X"7C", X"00", --0C18
  X"00", X"42", X"00", X"42", X"42", X"42", X"4A", X"00", --0C20
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0C28
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0C30
  X"00", X"00", X"08", X"3E", X"42", X"48", X"00", X"00", --0C38
  X"00", X"10", X"00", X"40", X"40", X"40", X"10", X"00", --0C40
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0C48
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0C50
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0C58
  X"00", X"18", X"00", X"7C", X"08", X"4E", X"42", X"10", --0C60
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0C68
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0C70
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0C78
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0C80
  X"00", X"00", X"00", X"02", X"40", X"42", X"7C", X"40", --0C88
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0C90
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0C98
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0CA0
  X"00", X"00", X"00", X"42", X"08", X"4E", X"42", X"00", --0CA8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0CB0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0CB8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0CC0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0CC8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0CD0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0CD8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0CE0
  X"00", X"00", X"02", X"7C", X"7E", X"40", X"40", X"00", --0CE8
  X"10", X"42", X"00", X"02", X"10", X"7E", X"7C", X"10", --0CF0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0CF8
  X"00", X"46", X"00", X"42", X"40", X"00", X"00", X"00", --0D00
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0D08
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"99", --0D10
  X"00", X"42", X"42", X"40", X"40", X"42", X"44", X"00", --0D18
  X"00", X"42", X"00", X"44", X"42", X"5A", X"46", X"00", --0D20
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0D28
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0D30
  X"00", X"00", X"08", X"02", X"42", X"7E", X"00", X"00", --0D38
  X"00", X"20", X"00", X"40", X"40", X"40", X"10", X"00", --0D40
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0D48
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0D50
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0D58
  X"00", X"24", X"00", X"44", X"08", X"42", X"42", X"10", --0D60
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0D68
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0D70
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0D78
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0D80
  X"00", X"00", X"00", X"42", X"42", X"42", X"44", X"40", --0D88
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0D90
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0D98
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0DA0
  X"00", X"00", X"00", X"42", X"08", X"42", X"42", X"00", --0DA8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0DB0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0DB8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0DC0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0DC8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0DD0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0DD8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0DE0
  X"00", X"00", X"42", X"40", X"42", X"42", X"40", X"00", --0DE8
  X"10", X"42", X"00", X"42", X"10", X"42", X"44", X"10", --0DF0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0DF8
  X"00", X"42", X"00", X"3C", X"40", X"00", X"00", X"00", --0E00
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0E08
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"42", --0E10
  X"00", X"7C", X"3C", X"7E", X"7E", X"42", X"42", X"00", --0E18
  X"00", X"42", X"00", X"78", X"3C", X"24", X"42", X"00", --0E20
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0E28
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0E30
  X"00", X"00", X"3E", X"3C", X"3C", X"08", X"00", X"00", --0E38
  X"00", X"7E", X"00", X"7E", X"7E", X"40", X"10", X"00", --0E40
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0E48
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0E50
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0E58
  X"00", X"42", X"00", X"42", X"3E", X"3C", X"42", X"10", --0E60
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0E68
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0E70
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0E78
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0E80
  X"00", X"00", X"00", X"3C", X"3C", X"3C", X"42", X"7E", --0E88
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0E90
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0E98
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0EA0
  X"00", X"00", X"00", X"42", X"3E", X"3C", X"42", X"00", --0EA8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0EB0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0EB8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0EC0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0EC8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0ED0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0ED8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0EE0
  X"00", X"00", X"3C", X"40", X"42", X"3C", X"7E", X"00", --0EE8
  X"10", X"3C", X"00", X"3C", X"10", X"42", X"42", X"10", --0EF0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0EF8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F00
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F08
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"3C", --0F10
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F18
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F20
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F28
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F30
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F38
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F40
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F48
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F50
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F58
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F60
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F68
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F70
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F78
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F80
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F88
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F90
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0F98
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0FA0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0FA8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0FB0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0FB8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0FC0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0FC8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0FD0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0FD8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0FE0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0FE8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0FF0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --0FF8
  X"00", X"3F", X"C0", X"00", X"00", X"00", X"00", X"00", --1000
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1008
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1010
  X"00", X"7C", X"00", X"00", X"00", X"FF", X"E0", X"00", --1018
  X"FF", X"FF", X"FF", X"80", X"00", X"00", X"60", X"04", --1020
  X"60", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1028
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1030
  X"3E", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1038
  X"FF", X"FF", X"FE", X"00", X"00", X"01", X"00", X"10", --1040
  X"00", X"00", X"00", X"00", X"3F", X"00", X"00", X"00", --1048
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1050
  X"3E", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1058
  X"FF", X"FF", X"FE", X"00", X"00", X"00", X"00", X"00", --1060
  X"00", X"00", X"00", X"00", X"FE", X"00", X"00", X"00", --1068
  X"00", X"3F", X"FF", X"FC", X"00", X"00", X"00", X"00", --1070
  X"7E", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1078
  X"FF", X"FF", X"FE", X"00", X"00", X"00", X"00", X"00", --1080
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1088
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1090
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1098
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --10A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --10A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --10B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --10B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --10C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --10C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --10D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --10D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --10E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --10E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --10F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --10F8
  X"00", X"FF", X"F0", X"00", X"00", X"00", X"00", X"00", --1100
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1108
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1110
  X"01", X"FF", X"00", X"00", X"03", X"FF", X"F8", X"00", --1118
  X"FF", X"FF", X"FF", X"F0", X"00", X"00", X"40", X"04", --1120
  X"F0", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1128
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1130
  X"3E", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1138
  X"FF", X"FF", X"FC", X"00", X"00", X"01", X"00", X"10", --1140
  X"00", X"00", X"00", X"00", X"3F", X"00", X"00", X"00", --1148
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1150
  X"1E", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1158
  X"FF", X"FF", X"FF", X"00", X"00", X"00", X"00", X"00", --1160
  X"00", X"00", X"00", X"00", X"FF", X"00", X"07", X"FF", --1168
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"E0", X"00", --1170
  X"FE", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1178
  X"FF", X"FF", X"FE", X"00", X"00", X"00", X"00", X"00", --1180
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1188
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1190
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1198
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --11A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --11A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --11B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --11B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --11C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --11C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --11D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --11D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --11E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --11E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --11F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --11F8
  X"3F", X"FF", X"F0", X"00", X"00", X"00", X"00", X"00", --1200
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1208
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1210
  X"07", X"FF", X"E0", X"00", X"0F", X"FF", X"FE", X"03", --1218
  X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"40", X"08", --1220
  X"F0", X"00", X"0F", X"FF", X"E0", X"00", X"00", X"00", --1228
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1230
  X"3E", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1238
  X"FF", X"FF", X"FC", X"00", X"00", X"01", X"00", X"10", --1240
  X"00", X"00", X"00", X"00", X"7F", X"00", X"00", X"00", --1248
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1250
  X"1E", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1258
  X"FF", X"FF", X"FF", X"00", X"00", X"00", X"00", X"00", --1260
  X"00", X"00", X"00", X"00", X"7F", X"FF", X"FF", X"FF", --1268
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1270
  X"FE", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1278
  X"FF", X"FF", X"FE", X"00", X"00", X"00", X"00", X"00", --1280
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1288
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1290
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1298
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --12A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --12A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --12B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --12B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --12C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --12C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --12D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --12D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --12E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --12E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --12F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --12F8
  X"FF", X"FF", X"F8", X"00", X"00", X"00", X"00", X"00", --1300
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1308
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1310
  X"1F", X"FF", X"F8", X"00", X"3F", X"FF", X"FF", X"FF", --1318
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"C0", X"08", --1320
  X"F0", X"03", X"FF", X"FF", X"F0", X"00", X"00", X"00", --1328
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1330
  X"7E", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1338
  X"FF", X"FF", X"FC", X"00", X"00", X"01", X"00", X"10", --1340
  X"00", X"00", X"00", X"00", X"7F", X"00", X"00", X"00", --1348
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1350
  X"1F", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1358
  X"FF", X"FF", X"FF", X"00", X"00", X"00", X"00", X"00", --1360
  X"00", X"00", X"00", X"00", X"3F", X"FF", X"FF", X"FF", --1368
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1370
  X"FC", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1378
  X"FF", X"FF", X"FC", X"00", X"00", X"00", X"00", X"00", --1380
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1388
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1390
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1398
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --13A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --13A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --13B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --13B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --13C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --13C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --13D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --13D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --13E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --13E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --13F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --13F8
  X"FF", X"FF", X"F8", X"00", X"00", X"00", X"0A", X"00", --1400
  X"60", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1408
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1410
  X"1F", X"FF", X"FF", X"FF", X"FF", X"E0", X"3F", X"FF", --1418
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"80", X"08", --1420
  X"FF", X"FF", X"FF", X"FF", X"FC", X"00", X"00", X"00", --1428
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1430
  X"7E", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1438
  X"FF", X"FF", X"FE", X"00", X"00", X"01", X"00", X"10", --1440
  X"00", X"00", X"00", X"00", X"7F", X"00", X"00", X"00", --1448
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1450
  X"1F", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1458
  X"FF", X"FF", X"FF", X"00", X"00", X"00", X"00", X"00", --1460
  X"00", X"00", X"00", X"00", X"3F", X"FF", X"FF", X"FF", --1468
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --1470
  X"F8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1478
  X"FF", X"FF", X"FC", X"00", X"00", X"00", X"00", X"00", --1480
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1488
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1490
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1498
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --14A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --14A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --14B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --14B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --14C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --14C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --14D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --14D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --14E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --14E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --14F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --14F8
  X"FF", X"FF", X"FC", X"00", X"00", X"00", X"10", X"01", --1500
  X"98", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1508
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1510
  X"3F", X"FF", X"FF", X"FF", X"FE", X"00", X"07", X"FE", --1518
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"80", X"08", --1520
  X"FF", X"FF", X"FF", X"FF", X"FE", X"00", X"00", X"00", --1528
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1530
  X"3E", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1538
  X"FF", X"FF", X"FE", X"00", X"00", X"00", X"00", X"00", --1540
  X"00", X"00", X"00", X"00", X"FE", X"00", X"00", X"00", --1548
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1550
  X"1F", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1558
  X"FF", X"FF", X"FF", X"00", X"00", X"00", X"00", X"00", --1560
  X"00", X"00", X"00", X"00", X"1F", X"FF", X"FF", X"FF", --1568
  X"FF", X"80", X"00", X"03", X"FF", X"FF", X"FF", X"FF", --1570
  X"F0", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1578
  X"FF", X"FF", X"FC", X"00", X"00", X"00", X"00", X"00", --1580
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1588
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1590
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1598
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --15A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --15A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --15B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --15B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --15C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --15C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --15D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --15D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --15E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --15E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --15F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --15F8
  X"FF", X"FF", X"FC", X"00", X"00", X"00", X"20", X"02", --1600
  X"04", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1608
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1610
  X"3F", X"C1", X"FF", X"FF", X"F0", X"00", X"00", X"FC", --1618
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"80", X"08", --1620
  X"FF", X"FF", X"FF", X"3F", X"FE", X"00", X"00", X"00", --1628
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1630
  X"3E", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1638
  X"FF", X"FF", X"FE", X"00", X"00", X"00", X"00", X"00", --1640
  X"00", X"00", X"00", X"00", X"FE", X"00", X"00", X"00", --1648
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1650
  X"3F", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1658
  X"FF", X"FF", X"FE", X"00", X"00", X"00", X"00", X"00", --1660
  X"00", X"00", X"00", X"00", X"07", X"FF", X"FF", X"C0", --1668
  X"00", X"00", X"00", X"00", X"00", X"03", X"FF", X"FF", --1670
  X"E0", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1678
  X"FF", X"FF", X"FC", X"00", X"00", X"00", X"00", X"00", --1680
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1688
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1690
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1698
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --16A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --16A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --16B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --16B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --16C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --16C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --16D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --16D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --16E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --16E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --16F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --16F8
  X"FF", X"FF", X"FF", X"00", X"00", X"00", X"20", X"04", --1700
  X"02", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1708
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1710
  X"3F", X"80", X"3F", X"FF", X"80", X"00", X"00", X"00", --1718
  X"FF", X"FF", X"FF", X"00", X"07", X"FC", X"80", X"08", --1720
  X"FF", X"FF", X"00", X"00", X"7F", X"00", X"00", X"00", --1728
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1730
  X"3E", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1738
  X"FF", X"FF", X"FE", X"00", X"00", X"00", X"00", X"00", --1740
  X"00", X"00", X"00", X"00", X"FE", X"00", X"00", X"00", --1748
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1750
  X"3F", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1758
  X"FF", X"FF", X"FE", X"00", X"00", X"00", X"00", X"00", --1760
  X"00", X"00", X"00", X"00", X"03", X"FF", X"00", X"00", --1768
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"FF", --1770
  X"C0", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1778
  X"FF", X"FF", X"FC", X"00", X"00", X"00", X"00", X"00", --1780
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1788
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1790
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1798
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --17A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --17A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --17B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --17B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --17C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --17C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --17D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --17D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --17E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --17E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --17F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --17F8
  X"00", X"00", X"36", X"00", X"36", X"00", X"36", X"00", --1800
  X"36", X"36", X"36", X"36", X"36", X"00", X"36", X"00", --1808
  X"00", X"00", X"00", X"36", X"36", X"36", X"36", X"00", --1810
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1818
  X"00", X"00", X"36", X"00", X"36", X"00", X"36", X"00", --1820
  X"36", X"00", X"00", X"00", X"36", X"00", X"36", X"00", --1828
  X"00", X"00", X"00", X"36", X"00", X"00", X"00", X"00", --1830
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1838
  X"00", X"00", X"36", X"00", X"36", X"00", X"36", X"00", --1840
  X"36", X"00", X"00", X"00", X"36", X"00", X"36", X"00", --1848
  X"00", X"00", X"00", X"36", X"36", X"36", X"00", X"00", --1850
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1858
  X"00", X"00", X"36", X"36", X"36", X"36", X"36", X"00", --1860
  X"36", X"36", X"36", X"36", X"36", X"00", X"36", X"36", --1868
  X"36", X"36", X"00", X"36", X"00", X"00", X"00", X"00", --1870
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1878
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1880
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1888
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1890
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1898
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --18A0
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --18A8
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --18B0
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --18B8
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --18C0
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --18C8
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --18D0
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --18D8
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --18E0
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --18E8
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --18F0
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --18F8
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1900
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1908
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1910
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1918
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1920
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1928
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1930
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1938
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1940
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1948
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1950
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1958
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1960
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1968
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1970
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1978
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1980
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1988
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1990
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --1998
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --19A0
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --19A8
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --19B0
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --19B8
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --19C0
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --19C8
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --19D0
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --19D8
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --19E0
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --19E8
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"42", --19F0
  X"42", X"42", X"42", X"42", X"42", X"42", X"42", X"00", --19F8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A00
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A08
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A10
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A18
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A20
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A28
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A30
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A38
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A40
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A48
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A50
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A58
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A60
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A68
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A70
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A78
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A80
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A88
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A90
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1A98
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1AA0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1AA8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1AB0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1AB8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1AC0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1AC8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1AD0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1AD8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1AE0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1AE8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1AF0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1AF8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B00
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B08
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B10
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B18
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B20
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B28
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B30
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B38
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B40
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B48
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B50
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B58
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B60
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B68
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B70
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B78
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B80
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B88
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B90
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1B98
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1BA0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1BA8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1BB0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1BB8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1BC0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1BC8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1BD0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1BD8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1BE0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1BE8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1BF0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1BF8
  X"FF", X"00", X"00", X"00", X"FF", X"00", X"23", X"0D", --1C00
  X"0D", X"23", X"05", X"00", X"00", X"00", X"10", X"0A", --1C08
  X"01", X"00", X"06", X"00", X"0B", X"00", X"01", X"00", --1C10
  X"01", X"00", X"06", X"00", X"10", X"00", X"00", X"00", --1C18
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1C20
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1C28
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"3C", --1C30
  X"40", X"00", X"FF", X"CD", X"00", X"20", X"5E", X"00", --1C38
  X"00", X"00", X"0A", X"00", X"FF", X"28", X"00", X"01", --1C40
  X"00", X"00", X"00", X"63", X"5D", X"00", X"00", X"B6", --1C48
  X"5C", X"BB", X"5C", X"CB", X"5C", X"63", X"5D", X"CA", --1C50
  X"5C", X"64", X"5D", X"67", X"5D", X"62", X"5D", X"BE", --1C58
  X"5D", X"69", X"5D", X"69", X"5D", X"69", X"5D", X"2D", --1C60
  X"92", X"5C", X"00", X"02", X"00", X"00", X"00", X"00", --1C68
  X"00", X"00", X"00", X"00", X"B6", X"1A", X"00", X"00", --1C70
  X"38", X"03", X"00", X"58", X"7F", X"00", X"00", X"21", --1C78
  X"00", X"5B", X"21", X"17", X"E0", X"48", X"E0", X"50", --1C80
  X"21", X"09", X"21", X"17", X"03", X"00", X"00", X"00", --1C88
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1C90
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1C98
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1CA0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1CA8
  X"00", X"00", X"23", X"5E", X"FF", X"7F", X"F4", X"09", --1CB0
  X"A8", X"10", X"4B", X"F4", X"09", X"C4", X"15", X"53", --1CB8
  X"81", X"0F", X"C4", X"15", X"52", X"F4", X"09", X"C4", --1CC0
  X"15", X"50", X"80", X"00", X"0A", X"0D", X"00", X"FD", --1CC8
  X"32", X"34", X"30", X"39", X"39", X"0E", X"00", X"00", --1CD0
  X"23", X"5E", X"00", X"0D", X"00", X"0B", X"09", X"00", --1CD8
  X"E7", X"30", X"0E", X"00", X"00", X"00", X"00", X"00", --1CE0
  X"0D", X"00", X"0F", X"14", X"00", X"D9", X"30", X"0E", --1CE8
  X"00", X"00", X"00", X"00", X"00", X"3A", X"DA", X"30", --1CF0
  X"0E", X"00", X"00", X"00", X"00", X"00", X"3A", X"FB", --1CF8
  X"0D", X"00", X"11", X"24", X"00", X"F5", X"AC", X"31", --1D00
  X"30", X"0E", X"00", X"00", X"0A", X"00", X"00", X"2C", --1D08
  X"31", X"30", X"0E", X"00", X"00", X"0A", X"00", X"00", --1D10
  X"3B", X"22", X"10", X"06", X"50", X"6C", X"65", X"61", --1D18
  X"73", X"65", X"20", X"57", X"61", X"69", X"74", X"22", --1D20
  X"0D", X"00", X"14", X"10", X"00", X"EF", X"22", X"22", --1D28
  X"AF", X"32", X"34", X"31", X"30", X"30", X"0E", X"00", --1D30
  X"00", X"24", X"5E", X"00", X"0D", X"00", X"1E", X"10", --1D38
  X"00", X"EF", X"22", X"22", X"AF", X"31", X"36", X"33", --1D40
  X"38", X"34", X"0E", X"00", X"00", X"00", X"40", X"00", --1D48
  X"0D", X"00", X"28", X"0E", X"00", X"F9", X"C0", X"32", --1D50
  X"35", X"30", X"30", X"30", X"0E", X"00", X"00", X"A8", --1D58
  X"61", X"00", X"0D", X"80", X"EF", X"22", X"22", X"0D", --1D60
  X"80", X"00", X"00", X"A8", X"61", X"00", X"20", X"20", --1D68
  X"20", X"20", X"20", X"20", X"00", X"00", X"00", X"40", --1D70
  X"00", X"00", X"03", X"57", X"6F", X"6F", X"6C", X"75", --1D78
  X"66", X"32", X"20", X"20", X"20", X"00", X"18", X"00", --1D80
  X"80", X"00", X"80", X"00", X"00", X"00", X"40", X"00", --1D88
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1D90
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1D98
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1DA0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1DA8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1DB0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1DB8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1DC0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1DC8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1DD0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1DD8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1DE0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1DE8
  X"00", X"00", X"DB", X"02", X"4D", X"00", X"DB", X"02", --1DF0
  X"4D", X"00", X"05", X"3D", X"00", X"04", X"DB", X"02", --1DF8
  X"4D", X"00", X"08", X"3D", X"00", X"00", X"00", X"00", --1E00
  X"09", X"DF", X"EE", X"64", X"2B", X"2D", X"65", X"33", --1E08
  X"00", X"00", X"ED", X"10", X"0D", X"00", X"09", X"00", --1E10
  X"85", X"1C", X"10", X"1C", X"52", X"1B", X"76", X"1B", --1E18
  X"03", X"13", X"00", X"3E", X"49", X"64", X"64", X"64", --1E20
  X"49", X"49", X"49", X"64", X"49", X"49", X"49", X"64", --1E28
  X"49", X"64", X"64", X"64", X"49", X"49", X"49", X"64", --1E30
  X"49", X"49", X"49", X"64", X"49", X"64", X"49", X"64", --1E38
  X"64", X"64", X"49", X"64", X"64", X"49", X"64", X"64", --1E40
  X"49", X"64", X"64", X"64", X"49", X"64", X"49", X"64", --1E48
  X"49", X"64", X"64", X"64", X"49", X"64", X"49", X"64", --1E50
  X"49", X"64", X"64", X"64", X"49", X"64", X"49", X"64", --1E58
  X"64", X"49", X"64", X"64", X"64", X"64", X"64", X"64", --1E60
  X"49", X"64", X"64", X"64", X"49", X"64", X"49", X"64", --1E68
  X"49", X"64", X"64", X"64", X"49", X"64", X"49", X"64", --1E70
  X"49", X"64", X"64", X"64", X"49", X"64", X"49", X"64", --1E78
  X"64", X"64", X"64", X"64", X"64", X"64", X"64", X"64", --1E80
  X"49", X"49", X"49", X"64", X"49", X"49", X"49", X"64", --1E88
  X"49", X"64", X"64", X"64", X"49", X"49", X"49", X"64", --1E90
  X"49", X"49", X"49", X"64", X"49", X"49", X"49", X"64", --1E98
  X"64", X"64", X"64", X"64", X"64", X"64", X"64", X"64", --1EA0
  X"64", X"64", X"49", X"64", X"49", X"64", X"64", X"64", --1EA8
  X"49", X"64", X"64", X"64", X"49", X"64", X"49", X"64", --1EB0
  X"64", X"64", X"49", X"64", X"49", X"64", X"49", X"64", --1EB8
  X"64", X"64", X"64", X"64", X"64", X"49", X"64", X"64", --1EC0
  X"64", X"64", X"49", X"64", X"49", X"64", X"64", X"64", --1EC8
  X"49", X"64", X"64", X"64", X"49", X"64", X"49", X"64", --1ED0
  X"64", X"64", X"49", X"64", X"49", X"64", X"49", X"64", --1ED8
  X"64", X"49", X"64", X"64", X"49", X"64", X"64", X"64", --1EE0
  X"49", X"49", X"49", X"64", X"49", X"64", X"64", X"64", --1EE8
  X"49", X"49", X"49", X"64", X"49", X"64", X"49", X"64", --1EF0
  X"49", X"49", X"49", X"64", X"49", X"64", X"49", X"64", --1EF8
  X"64", X"64", X"49", X"64", X"64", X"64", X"64", X"64", --1F00
  X"64", X"64", X"64", X"64", X"64", X"64", X"64", X"64", --1F08
  X"64", X"64", X"64", X"64", X"64", X"64", X"64", X"64", --1F10
  X"64", X"64", X"64", X"64", X"64", X"64", X"64", X"64", --1F18
  X"64", X"64", X"64", X"4E", X"00", X"00", X"36", X"00", --1F20
  X"36", X"00", X"36", X"00", X"36", X"36", X"36", X"36", --1F28
  X"36", X"00", X"36", X"00", X"00", X"00", X"00", X"36", --1F30
  X"36", X"36", X"36", X"00", X"00", X"00", X"00", X"00", --1F38
  X"00", X"00", X"00", X"00", X"00", X"00", X"36", X"00", --1F40
  X"36", X"00", X"36", X"00", X"36", X"00", X"00", X"00", --1F48
  X"36", X"00", X"36", X"00", X"00", X"00", X"00", X"36", --1F50
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1F58
  X"00", X"00", X"00", X"00", X"00", X"00", X"36", X"00", --1F60
  X"36", X"00", X"36", X"00", X"36", X"00", X"00", X"00", --1F68
  X"36", X"00", X"36", X"00", X"00", X"00", X"00", X"36", --1F70
  X"36", X"36", X"00", X"00", X"00", X"00", X"00", X"00", --1F78
  X"00", X"00", X"00", X"00", X"00", X"00", X"36", X"36", --1F80
  X"36", X"36", X"36", X"00", X"36", X"36", X"36", X"36", --1F88
  X"36", X"00", X"36", X"36", X"36", X"36", X"00", X"36", --1F90
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1F98
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1FA0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1FA8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1FB0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --1FB8
  X"00", X"00", X"CE", X"0B", X"E5", X"50", X"CE", X"0B", --1FC0
  X"E6", X"50", X"1B", X"17", X"DC", X"0A", X"CE", X"0B", --1FC8
  X"E9", X"50", X"18", X"17", X"DC", X"0A", X"D7", X"18", --1FD0
  X"38", X"00", X"B1", X"33", X"15", X"5D", X"DB", X"02", --1FD8
  X"4D", X"00", X"84", X"4F", X"7C", X"00", X"83", X"4F", --1FE0
  X"8C", X"10", X"5C", X"0E", X"00", X"47", X"C0", X"57", --1FE8
  X"71", X"0E", X"F3", X"0D", X"21", X"17", X"C6", X"1E", --1FF0
  X"1A", X"5E", X"76", X"1B", X"03", X"13", X"00", X"3E", --1FF8
  X"C3", X"3A", X"61", X"16", X"75", X"DD", X"87", X"D4", --2000
  X"03", X"3A", X"5C", X"E8", X"5F", X"E1", X"A7", X"3E", --2008
  X"0D", X"3F", X"0D", X"45", X"4F", X"46", X"0D", X"4D", --2010
  X"45", X"4D", X"4F", X"52", X"59", X"0D", X"52", X"45", --2018
  X"53", X"45", X"52", X"56", X"45", X"44", X"0D", X"46", --2020
  X"55", X"4C", X"4C", X"0D", X"44", X"4F", X"55", X"42", --2028
  X"4C", X"45", X"0D", X"53", X"59", X"4D", X"42", X"4F", --2030
  X"4C", X"0D", X"4F", X"50", X"45", X"52", X"41", X"4E", --2038
  X"44", X"0D", X"55", X"4E", X"44", X"45", X"46", X"49", --2040
  X"4E", X"45", X"44", X"0D", X"4F", X"52", X"47", X"2D", --2048
  X"0D", X"2A", X"2A", X"2A", X"2A", X"2A", X"2A", X"2A", --2050
  X"2A", X"20", X"41", X"53", X"50", X"45", X"43", X"54", --2058
  X"20", X"34", X"2E", X"32", X"20", X"2A", X"2A", X"2A", --2060
  X"2A", X"2A", X"2A", X"2A", X"2A", X"0D", X"CB", X"F5", --2068
  X"CE", X"FE", X"55", X"20", X"04", X"DD", X"CB", X"F5", --2070
  X"E6", X"FE", X"41", X"20", X"E6", X"DD", X"CB", X"F5", --2078
  X"C6", X"1A", X"FE", X"20", X"20", X"03", X"13", X"18", --2080
  X"DB", X"02", X"4D", X"00", X"DB", X"02", X"DB", X"02", --2088
  X"DB", X"02", X"DB", X"02", X"4D", X"00", X"91", X"47", --2090
  X"DB", X"02", X"4D", X"00", X"8A", X"4E", X"56", X"00", --2098
  X"AA", X"4E", X"0D", X"0F", X"E0", X"57", X"71", X"0E", --20A0
  X"DF", X"0C", X"F3", X"0D", X"CE", X"0B", X"F3", X"0D", --20A8
  X"F3", X"0D", X"21", X"02", X"FE", X"15", X"58", X"27", --20B0
  X"8A", X"63", X"4E", X"63", X"16", X"61", X"4A", X"0D", --20B8
  X"CF", X"60", X"F4", X"60", X"02", X"00", X"71", X"63", --20C0
  X"4A", X"52", X"72", X"61", X"61", X"61", X"52", X"0D", --20C8
  X"30", X"0D", X"07", X"00", X"00", X"00", X"39", X"35", --20D0
  X"35", X"31", X"0D", X"35", X"0D", X"32", X"2C", X"30", --20D8
  X"2C", X"30", X"2C", X"30", X"0D", X"0D", X"2C", X"31", --20E0
  X"36", X"30", X"0D", X"32", X"0D", X"35", X"06", X"01", --20E8
  X"D9", X"3E", X"30", X"30", X"32", X"30", X"20", X"0D", --20F0
  X"0D", X"B7", X"20", X"53", X"21", X"22", X"12", X"CD", --20F8
  X"91", X"08", X"CD", X"BD", X"0B", X"7E", X"23", X"FE", --2100
  X"0D", X"28", X"1A", X"FE", X"41", X"20", X"04", X"DD", --2108
  X"CB", X"F5", X"C6", X"FE", X"43", X"20", X"56", X"09", --2110
  X"00", X"01", X"03", X"00", X"1F", X"08", X"05", X"06", --2118
  X"05", X"05", X"08", X"05", X"00", X"00", X"14", X"00", --2120
  X"00", X"FF", X"CC", X"75", X"00", X"00", X"DC", X"87", --2128
  X"BD", X"70", X"CC", X"60", X"BC", X"70", X"60", X"7F", --2130
  X"E0", X"D6", X"DD", X"22", X"07", X"60", X"FD", X"22", --2138
  X"09", X"60", X"ED", X"73", X"0B", X"60", X"31", X"CE", --2140
  X"60", X"CD", X"BA", X"65", X"22", X"28", X"61", X"DD", --2148
  X"21", X"16", X"61", X"CD", X"E5", X"61", X"CD", X"6B", --2150
  X"63", X"2E", X"51", X"CD", X"ED", X"64", X"CD", X"6B", --2158
  X"63", X"21", X"61", X"61", X"E5", X"ED", X"73", X"32", --2160
  X"61", X"DD", X"36", X"00", X"56", X"2E", X"0F", X"CD", --2168
  X"F9", X"64", X"0D", X"C8", X"FE", X"53", X"CA", X"CF", --2170
  X"62", X"FE", X"48", X"CA", X"A7", X"61", X"FE", X"52", --2178
  X"CA", X"35", X"6F", X"E5", X"C5", X"0E", X"01", X"11", --2180
  X"CE", X"60", X"21", X"31", X"63", X"CD", X"72", X"68", --2188
  X"DA", X"56", X"65", X"C1", X"E3", X"41", X"05", X"37", --2190
  X"28", X"09", X"13", X"CD", X"5B", X"65", X"DA", X"56", --2198
  X"65", X"44", X"4D", X"2A", X"2A", X"61", X"C9", X"0D", --21A0
  X"C3", X"AF", X"64", X"00", X"00", X"B5", X"48", X"00", --21A8
  X"00", X"00", X"00", X"00", X"00", X"0A", X"00", X"00", --21B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --21B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --21C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --21C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"80", --21D0
  X"00", X"11", X"00", X"58", X"21", X"24", X"5F", X"ED", --21D8
  X"B0", X"C9", X"01", X"80", X"00", X"11", X"85", X"58", --21E0
  X"21", X"24", X"5F", X"7E", X"3C", X"3D", X"20", X"02", --21E8
  X"3E", X"64", X"CB", X"F7", X"12", X"23", X"13", X"0D", --21F0
  X"20", X"F1", X"C9", X"21", X"80", X"58", X"0E", X"80", --21F8
  X"3E", X"42", X"77", X"23", X"0D", X"20", X"FB", X"0E", --2200
  X"FF", X"77", X"23", X"0D", X"20", X"FB", X"3E", X"00", --2208
  X"0E", X"FF", X"77", X"23", X"0D", X"20", X"FB", X"77", --2210
  X"23", X"77", X"23", X"77", X"C9", X"21", X"70", X"59", --2218
  X"3E", X"64", X"77", X"ED", X"5B", X"B1", X"61", X"13", --2220
  X"ED", X"53", X"B1", X"61", X"21", X"00", X"58", X"01", --2228
  X"05", X"00", X"09", X"01", X"16", X"00", X"CD", X"45", --2230
  X"62", X"D5", X"11", X"21", X"00", X"19", X"D1", X"13", --2238
  X"0D", X"0D", X"20", X"F2", X"C9", X"C5", X"CD", X"5A", --2240
  X"62", X"C1", X"C5", X"CD", X"63", X"62", X"C1", X"C5", --2248
  X"CD", X"71", X"62", X"C1", X"C5", X"CD", X"7A", X"62", --2250
  X"C1", X"C9", X"1A", X"CB", X"BF", X"23", X"77", X"0D", --2258
  X"20", X"F8", X"C9", X"1A", X"CB", X"BF", X"D5", X"11", --2260
  X"20", X"00", X"19", X"D1", X"77", X"0D", X"20", X"F3", --2268
  X"C9", X"1A", X"CB", X"BF", X"2B", X"77", X"0D", X"20", --2270
  X"F8", X"C9", X"1A", X"CB", X"BF", X"D5", X"11", X"20", --2278
  X"00", X"ED", X"52", X"D1", X"77", X"0D", X"20", X"F2", --2280
  X"C9", X"00", X"49", X"52", X"5B", X"52", X"49", X"00", --2288
  X"49", X"52", X"5B", X"52", X"49", X"00", X"49", X"52", --2290
  X"5B", X"52", X"49", X"00", X"49", X"52", X"5B", X"52", --2298
  X"49", X"00", X"49", X"52", X"5B", X"52", X"49", X"00", --22A0
  X"49", X"52", X"5B", X"52", X"49", X"00", X"49", X"52", --22A8
  X"5B", X"52", X"49", X"00", X"49", X"52", X"5B", X"52", --22B0
  X"49", X"00", X"49", X"52", X"5B", X"52", X"49", X"00", --22B8
  X"49", X"52", X"5B", X"52", X"49", X"00", X"49", X"52", --22C0
  X"5B", X"52", X"49", X"00", X"49", X"52", X"5B", X"52", --22C8
  X"49", X"00", X"49", X"52", X"5B", X"52", X"49", X"00", --22D0
  X"49", X"52", X"5B", X"64", X"64", X"64", X"64", X"64", --22D8
  X"64", X"64", X"64", X"64", X"64", X"64", X"64", X"64", --22E0
  X"64", X"21", X"30", X"75", X"01", X"40", X"00", X"09", --22E8
  X"3E", X"67", X"0E", X"FF", X"77", X"23", X"0D", X"20", --22F0
  X"FB", X"0E", X"C1", X"77", X"23", X"0D", X"20", X"FB", --22F8
  X"01", X"C0", X"00", X"09", X"23", X"0E", X"40", X"77", --2300
  X"23", X"0D", X"20", X"FB", X"C9", X"21", X"40", X"40", --2308
  X"0E", X"06", X"C5", X"E5", X"CD", X"3B", X"63", X"E1", --2310
  X"01", X"20", X"00", X"09", X"C1", X"0D", X"20", X"F2", --2318
  X"21", X"80", X"42", X"CD", X"3B", X"63", X"21", X"A0", --2320
  X"42", X"CD", X"3B", X"63", X"21", X"C0", X"50", X"CD", --2328
  X"3B", X"63", X"21", X"E0", X"50", X"CD", X"3B", X"63", --2330
  X"C3", X"54", X"63", X"0E", X"08", X"C5", X"CD", X"4A", --2338
  X"63", X"01", X"E0", X"00", X"09", X"C1", X"0D", X"20", --2340
  X"F4", X"C9", X"0E", X"20", X"3E", X"00", X"77", X"23", --2348
  X"0D", X"20", X"F9", X"C9", X"21", X"00", X"48", X"0E", --2350
  X"08", X"C5", X"CD", X"62", X"63", X"C1", X"0D", X"20", --2358
  X"F8", X"C9", X"0E", X"FF", X"3E", X"00", X"77", X"23", --2360
  X"0D", X"20", X"F9", X"77", X"23", X"C9", X"21", X"31", --2368
  X"78", X"11", X"00", X"58", X"01", X"00", X"03", X"ED", --2370
  X"B0", X"21", X"00", X"58", X"01", X"0A", X"01", X"09", --2378
  X"3E", X"70", X"77", X"23", X"77", X"23", X"77", X"23", --2380
  X"77", X"01", X"05", X"00", X"09", X"77", X"23", X"77", --2388
  X"23", X"77", X"23", X"77", X"3E", X"56", X"CD", X"D3", --2390
  X"63", X"CD", X"11", X"64", X"CD", X"11", X"64", X"3E", --2398
  X"56", X"CD", X"D3", X"63", X"3E", X"62", X"CD", X"D3", --23A0
  X"63", X"CD", X"11", X"64", X"CD", X"11", X"64", X"3E", --23A8
  X"62", X"CD", X"D3", X"63", X"3E", X"5C", X"CD", X"D3", --23B0
  X"63", X"CD", X"11", X"64", X"CD", X"11", X"64", X"3E", --23B8
  X"12", X"CD", X"F4", X"63", X"CD", X"11", X"64", X"3E", --23C0
  X"70", X"CD", X"F4", X"63", X"CD", X"11", X"64", X"CD", --23C8
  X"11", X"64", X"C9", X"21", X"CB", X"61", X"77", X"21", --23D0
  X"CC", X"61", X"3E", X"7F", X"77", X"21", X"3E", X"6E", --23D8
  X"CD", X"83", X"6D", X"21", X"CB", X"61", X"7E", X"C6", --23E0
  X"40", X"77", X"21", X"3E", X"6E", X"22", X"C9", X"61", --23E8
  X"CD", X"83", X"6D", X"C9", X"21", X"00", X"58", X"01", --23F0
  X"EB", X"00", X"09", X"77", X"23", X"77", X"01", X"1E", --23F8
  X"00", X"09", X"77", X"23", X"77", X"23", X"77", X"23", --2400
  X"77", X"01", X"1E", X"00", X"09", X"77", X"23", X"77", --2408
  X"C9", X"21", X"DC", X"05", X"11", X"14", X"00", X"CD", --2410
  X"B5", X"03", X"21", X"D0", X"07", X"11", X"0D", X"00", --2418
  X"CD", X"B5", X"03", X"C9", X"21", X"90", X"48", X"22", --2420
  X"AD", X"61", X"18", X"14", X"2A", X"B6", X"61", X"22", --2428
  X"AF", X"61", X"21", X"B0", X"48", X"22", X"AD", X"61", --2430
  X"18", X"06", X"21", X"17", X"40", X"22", X"AD", X"61", --2438
  X"21", X"AB", X"61", X"CB", X"8E", X"2A", X"AF", X"61", --2440
  X"01", X"10", X"27", X"CD", X"67", X"64", X"01", X"E8", --2448
  X"03", X"CD", X"67", X"64", X"01", X"64", X"00", X"CD", --2450
  X"67", X"64", X"01", X"0A", X"00", X"CD", X"67", X"64", --2458
  X"01", X"01", X"00", X"CD", X"67", X"64", X"C9", X"AF", --2460
  X"ED", X"42", X"3C", X"30", X"FB", X"09", X"3D", X"20", --2468
  X"0F", X"3A", X"AB", X"61", X"CB", X"4F", X"20", X"04", --2470
  X"3E", X"20", X"18", X"0D", X"3E", X"4F", X"18", X"09", --2478
  X"E5", X"21", X"AB", X"61", X"CB", X"CE", X"E1", X"C6", --2480
  X"30", X"E5", X"CD", X"99", X"64", X"21", X"AD", X"61", --2488
  X"34", X"2A", X"AD", X"61", X"CD", X"A6", X"64", X"E1", --2490
  X"C9", X"ED", X"4B", X"36", X"5C", X"26", X"00", X"6F", --2498
  X"29", X"29", X"29", X"09", X"EB", X"C9", X"06", X"08", --24A0
  X"1A", X"77", X"24", X"13", X"10", X"FA", X"C9", X"21", --24A8
  X"48", X"5C", X"3E", X"00", X"77", X"21", X"00", X"00", --24B0
  X"22", X"B6", X"61", X"22", X"AF", X"61", X"21", X"B5", --24B8
  X"61", X"3E", X"0A", X"77", X"3E", X"00", X"0E", X"FE", --24C0
  X"ED", X"79", X"CD", X"D6", X"61", X"CD", X"FB", X"61", --24C8
  X"CD", X"0D", X"63", X"CD", X"EA", X"65", X"CD", X"24", --24D0
  X"64", X"2A", X"AF", X"61", X"ED", X"4B", X"B6", X"61", --24D8
  X"AF", X"ED", X"42", X"38", X"06", X"2A", X"AF", X"61", --24E0
  X"22", X"B6", X"61", X"CD", X"2C", X"64", X"3E", X"7F", --24E8
  X"DB", X"FE", X"1F", X"DA", X"EE", X"64", X"21", X"70", --24F0
  X"73", X"3E", X"00", X"77", X"CD", X"0D", X"63", X"CD", --24F8
  X"6E", X"63", X"CD", X"0D", X"63", X"21", X"89", X"62", --2500
  X"22", X"B1", X"61", X"0E", X"53", X"C5", X"CD", X"CD", --2508
  X"6A", X"CD", X"1D", X"62", X"11", X"14", X"00", X"C1", --2510
  X"C5", X"26", X"01", X"79", X"C6", X"32", X"6F", X"CD", --2518
  X"B5", X"03", X"C1", X"0D", X"20", X"E7", X"21", X"AF", --2520
  X"61", X"11", X"00", X"00", X"ED", X"53", X"AF", X"61", --2528
  X"CD", X"3A", X"64", X"21", X"01", X"58", X"22", X"B8", --2530
  X"61", X"21", X"B3", X"61", X"3E", X"FF", X"77", X"21", --2538
  X"B4", X"61", X"3E", X"AF", X"77", X"21", X"AB", X"61", --2540
  X"CB", X"C6", X"CB", X"BE", X"CD", X"0D", X"63", X"21", --2548
  X"70", X"73", X"34", X"7E", X"D6", X"04", X"21", X"C3", --2550
  X"61", X"20", X"04", X"3E", X"08", X"18", X"03", X"3A", --2558
  X"B5", X"61", X"77", X"3E", X"00", X"21", X"B5", X"61", --2560
  X"77", X"CD", X"E9", X"62", X"CD", X"C1", X"6A", X"CD", --2568
  X"32", X"6B", X"CD", X"B7", X"6A", X"CD", X"E6", X"6C", --2570
  X"CD", X"C1", X"6A", X"CD", X"A5", X"6C", X"CD", X"4C", --2578
  X"6C", X"CD", X"0B", X"66", X"CD", X"90", X"6F", X"CD", --2580
  X"5A", X"71", X"CD", X"72", X"7B", X"21", X"AB", X"61", --2588
  X"CB", X"46", X"28", X"1A", X"CB", X"86", X"21", X"AB", --2590
  X"61", X"CB", X"7E", X"28", X"03", X"CD", X"CD", X"65", --2598
  X"CD", X"8E", X"6F", X"CD", X"09", X"66", X"CD", X"CD", --25A0
  X"65", X"CD", X"8E", X"6F", X"18", X"DF", X"CD", X"CD", --25A8
  X"6A", X"CD", X"8F", X"70", X"CD", X"E2", X"61", X"0E", --25B0
  X"14", X"CD", X"CD", X"6A", X"0D", X"20", X"FA", X"CD", --25B8
  X"10", X"72", X"21", X"AB", X"61", X"CB", X"7E", X"C2", --25C0
  X"39", X"65", X"C3", X"BE", X"64", X"CD", X"A3", X"69", --25C8
  X"21", X"71", X"73", X"77", X"CD", X"70", X"7B", X"21", --25D0
  X"72", X"73", X"CB", X"4E", X"28", X"0B", X"CD", X"C1", --25D8
  X"6A", X"CD", X"5A", X"71", X"21", X"72", X"73", X"CB", --25E0
  X"8E", X"C9", X"21", X"38", X"6F", X"7E", X"3C", X"3D", --25E8
  X"C8", X"23", X"3D", X"20", X"0C", X"7E", X"23", X"11", --25F0
  X"AD", X"61", X"12", X"13", X"7E", X"12", X"23", X"18", --25F8
  X"EC", X"3C", X"E5", X"CD", X"89", X"64", X"E1", X"18", --2600
  X"E4", X"18", X"2F", X"21", X"C4", X"61", X"3A", X"C3", --2608
  X"61", X"77", X"21", X"22", X"73", X"E5", X"E1", X"7E", --2610
  X"11", X"CB", X"61", X"12", X"23", X"7E", X"11", X"CC", --2618
  X"61", X"12", X"23", X"E5", X"01", X"D8", X"74", X"CD", --2620
  X"97", X"68", X"E1", X"3A", X"C9", X"61", X"77", X"23", --2628
  X"23", X"E5", X"21", X"C4", X"61", X"35", X"20", X"DE", --2630
  X"E1", X"C9", X"21", X"C4", X"61", X"3A", X"C3", X"61", --2638
  X"77", X"21", X"22", X"73", X"E5", X"E1", X"22", X"BF", --2640
  X"61", X"11", X"CB", X"61", X"7E", X"12", X"11", X"C7", --2648
  X"61", X"12", X"23", X"11", X"CC", X"61", X"7E", X"12", --2650
  X"11", X"C8", X"61", X"12", X"23", X"11", X"C9", X"61", --2658
  X"7E", X"12", X"11", X"C5", X"61", X"12", X"23", X"11", --2660
  X"C0", X"61", X"7E", X"12", X"E5", X"3A", X"C0", X"61", --2668
  X"CB", X"7F", X"20", X"03", X"CD", X"98", X"66", X"E1", --2670
  X"2B", X"2B", X"2B", X"3A", X"CB", X"61", X"77", X"23", --2678
  X"3A", X"CC", X"61", X"77", X"23", X"3A", X"C9", X"61", --2680
  X"77", X"23", X"3A", X"C0", X"61", X"77", X"23", X"E5", --2688
  X"21", X"C4", X"61", X"35", X"20", X"AF", X"E1", X"C9", --2690
  X"3A", X"C3", X"61", X"21", X"BE", X"61", X"77", X"21", --2698
  X"22", X"73", X"CD", X"A3", X"69", X"D6", X"0A", X"DA", --26A0
  X"9C", X"67", X"3A", X"BF", X"61", X"95", X"CA", X"9C", --26A8
  X"67", X"3A", X"CB", X"61", X"4F", X"7E", X"91", X"4F", --26B0
  X"23", X"3A", X"CC", X"61", X"47", X"7E", X"23", X"23", --26B8
  X"CB", X"7E", X"C2", X"9C", X"67", X"E5", X"21", X"C0", --26C0
  X"61", X"90", X"47", X"ED", X"43", X"C1", X"61", X"3A", --26C8
  X"C1", X"61", X"D6", X"1E", X"38", X"05", X"D6", X"C2", --26D0
  X"DA", X"9B", X"67", X"3A", X"C2", X"61", X"D6", X"1E", --26D8
  X"38", X"05", X"D6", X"C2", X"DA", X"9B", X"67", X"3A", --26E0
  X"C1", X"61", X"D6", X"0A", X"38", X"04", X"D6", X"EA", --26E8
  X"38", X"5F", X"3A", X"C2", X"61", X"D6", X"08", X"38", --26F0
  X"04", X"D6", X"EE", X"38", X"54", X"11", X"BE", X"61", --26F8
  X"3E", X"01", X"12", X"11", X"BE", X"61", X"3E", X"01", --2700
  X"12", X"3A", X"C1", X"61", X"D6", X"05", X"30", X"04", --2708
  X"CB", X"E6", X"18", X"19", X"D6", X"F5", X"38", X"04", --2710
  X"CB", X"E6", X"18", X"11", X"3A", X"C2", X"61", X"D6", --2718
  X"04", X"30", X"04", X"CB", X"E6", X"18", X"06", X"D6", --2720
  X"F7", X"38", X"02", X"CB", X"E6", X"3A", X"C1", X"61", --2728
  X"D6", X"0A", X"30", X"06", X"CB", X"8E", X"CB", X"C6", --2730
  X"18", X"04", X"CB", X"CE", X"CB", X"86", X"3A", X"C2", --2738
  X"61", X"D6", X"08", X"30", X"06", X"CB", X"96", X"CB", --2740
  X"DE", X"18", X"50", X"CB", X"9E", X"CB", X"D6", X"18", --2748
  X"4A", X"3A", X"C1", X"61", X"D6", X"0A", X"30", X"06", --2750
  X"CB", X"86", X"CB", X"8E", X"18", X"18", X"D6", X"14", --2758
  X"30", X"06", X"CB", X"CE", X"CB", X"86", X"18", X"0E", --2760
  X"D6", X"D6", X"30", X"06", X"CB", X"C6", X"CB", X"8E", --2768
  X"18", X"04", X"CB", X"86", X"CB", X"8E", X"3A", X"C2", --2770
  X"61", X"D6", X"08", X"30", X"06", X"CB", X"9E", X"CB", --2778
  X"96", X"18", X"18", X"D6", X"16", X"30", X"06", X"CB", --2780
  X"D6", X"CB", X"9E", X"18", X"0E", X"D6", X"D8", X"30", --2788
  X"06", X"CB", X"DE", X"CB", X"96", X"18", X"04", X"CB", --2790
  X"9E", X"CB", X"96", X"E1", X"23", X"E5", X"21", X"BE", --2798
  X"61", X"35", X"E1", X"C2", X"A2", X"66", X"CD", X"AB", --27A0
  X"6B", X"CB", X"50", X"28", X"13", X"CD", X"A3", X"69", --27A8
  X"D6", X"32", X"30", X"0F", X"CD", X"B9", X"69", X"21", --27B0
  X"C0", X"61", X"CB", X"AE", X"CB", X"A6", X"18", X"03", --27B8
  X"CD", X"B9", X"69", X"CD", X"86", X"6E", X"CD", X"DA", --27C0
  X"67", X"CD", X"3E", X"6B", X"CD", X"11", X"6F", X"CD", --27C8
  X"88", X"6A", X"21", X"C0", X"61", X"CB", X"7E", X"C0", --27D0
  X"18", X"1B", X"CD", X"A3", X"69", X"D6", X"03", X"30", --27D8
  X"13", X"CD", X"A3", X"69", X"E6", X"0F", X"21", X"C0", --27E0
  X"61", X"77", X"CB", X"46", X"28", X"06", X"CB", X"4E", --27E8
  X"28", X"02", X"18", X"E6", X"C9", X"21", X"AB", X"61", --27F0
  X"CB", X"C6", X"21", X"C0", X"61", X"CB", X"5E", X"28", --27F8
  X"13", X"3A", X"CC", X"61", X"D6", X"0C", X"30", X"06", --2800
  X"CB", X"9E", X"CB", X"D6", X"18", X"C4", X"21", X"CC", --2808
  X"61", X"35", X"18", X"18", X"21", X"C0", X"61", X"CB", --2810
  X"56", X"28", X"11", X"3A", X"CC", X"61", X"D6", X"AE", --2818
  X"38", X"06", X"CB", X"96", X"CB", X"DE", X"18", X"AA", --2820
  X"21", X"CC", X"61", X"34", X"21", X"C0", X"61", X"CB", --2828
  X"4E", X"28", X"15", X"3A", X"CB", X"61", X"D6", X"EE", --2830
  X"DA", X"42", X"68", X"CB", X"8E", X"CB", X"C6", X"C3", --2838
  X"D2", X"67", X"21", X"CB", X"61", X"34", X"18", X"19", --2840
  X"21", X"C0", X"61", X"CB", X"46", X"28", X"12", X"3A", --2848
  X"CB", X"61", X"D6", X"02", X"30", X"07", X"CB", X"86", --2850
  X"CB", X"CE", X"C3", X"D2", X"67", X"21", X"CB", X"61", --2858
  X"35", X"21", X"C0", X"61", X"CB", X"66", X"CB", X"A6", --2860
  X"C2", X"F5", X"67", X"CB", X"6E", X"CB", X"AE", X"C2", --2868
  X"F5", X"67", X"21", X"C9", X"61", X"3A", X"CB", X"61", --2870
  X"4F", X"3A", X"C7", X"61", X"91", X"28", X"0C", X"30", --2878
  X"04", X"CB", X"DE", X"18", X"02", X"CB", X"9E", X"CD", --2880
  X"C6", X"68", X"C9", X"3A", X"CC", X"61", X"4F", X"3A", --2888
  X"C8", X"61", X"91", X"28", X"F5", X"18", X"F0", X"ED", --2890
  X"43", X"C9", X"61", X"ED", X"43", X"C5", X"61", X"2A", --2898
  X"CB", X"61", X"22", X"C7", X"61", X"CD", X"16", X"69", --28A0
  X"C9", X"2A", X"CB", X"61", X"ED", X"4B", X"C7", X"61", --28A8
  X"ED", X"43", X"CB", X"61", X"22", X"C7", X"61", X"2A", --28B0
  X"C9", X"61", X"ED", X"4B", X"C5", X"61", X"22", X"C5", --28B8
  X"61", X"ED", X"43", X"C9", X"61", X"C9", X"CD", X"D2", --28C0
  X"68", X"ED", X"4B", X"CB", X"61", X"ED", X"43", X"C7", --28C8
  X"61", X"C9", X"2A", X"C9", X"61", X"E5", X"2A", X"CC", --28D0
  X"61", X"E5", X"2A", X"C5", X"61", X"E5", X"2A", X"C8", --28D8
  X"61", X"E5", X"0E", X"06", X"C5", X"CD", X"39", X"69", --28E0
  X"21", X"C9", X"61", X"34", X"21", X"CC", X"61", X"35", --28E8
  X"CD", X"A9", X"68", X"CD", X"39", X"69", X"21", X"C9", --28F0
  X"61", X"34", X"21", X"CC", X"61", X"35", X"CD", X"A9", --28F8
  X"68", X"C1", X"0D", X"20", X"DF", X"E1", X"22", X"C8", --2900
  X"61", X"E1", X"22", X"C5", X"61", X"E1", X"22", X"CC", --2908
  X"61", X"E1", X"22", X"C9", X"61", X"C9", X"2A", X"C9", --2910
  X"61", X"E5", X"2A", X"CC", X"61", X"E5", X"0E", X"06", --2918
  X"C5", X"CD", X"39", X"69", X"21", X"C9", X"61", X"34", --2920
  X"21", X"CC", X"61", X"35", X"C1", X"0D", X"20", X"F0", --2928
  X"E1", X"22", X"CC", X"61", X"E1", X"22", X"C9", X"61", --2930
  X"C9", X"3A", X"CC", X"61", X"C6", X"08", X"F5", X"0F", --2938
  X"0F", X"0F", X"E6", X"1F", X"47", X"3E", X"18", X"98", --2940
  X"47", X"3A", X"CB", X"61", X"0F", X"0F", X"0F", X"E6", --2948
  X"1F", X"4F", X"F1", X"E6", X"07", X"5F", X"3E", X"07", --2950
  X"9B", X"CD", X"90", X"69", X"3A", X"CB", X"61", X"E6", --2958
  X"07", X"4F", X"0C", X"0D", X"28", X"22", X"3E", X"FF", --2960
  X"C5", X"1F", X"CB", X"BF", X"0D", X"20", X"FA", X"57", --2968
  X"ED", X"4B", X"C9", X"61", X"0A", X"C1", X"0F", X"0D", --2970
  X"20", X"FC", X"5F", X"A2", X"AE", X"77", X"23", X"3E", --2978
  X"FF", X"AA", X"57", X"7B", X"A2", X"AE", X"77", X"C9", --2980
  X"ED", X"4B", X"C9", X"61", X"0A", X"AE", X"77", X"C9", --2988
  X"F5", X"78", X"E6", X"18", X"F6", X"40", X"67", X"F1", --2990
  X"84", X"67", X"78", X"E6", X"07", X"0F", X"0F", X"0F", --2998
  X"81", X"6F", X"C9", X"E5", X"21", X"BC", X"61", X"34", --29A0
  X"21", X"98", X"66", X"3A", X"BC", X"61", X"6F", X"3A", --29A8
  X"78", X"5C", X"86", X"21", X"79", X"5C", X"86", X"E1", --29B0
  X"C9", X"3A", X"CB", X"61", X"4F", X"3A", X"D5", X"61", --29B8
  X"91", X"4F", X"3A", X"CC", X"61", X"47", X"3A", X"D4", --29C0
  X"61", X"21", X"C0", X"61", X"90", X"47", X"ED", X"43", --29C8
  X"BA", X"61", X"3A", X"BA", X"61", X"D6", X"1E", X"38", --29D0
  X"05", X"D6", X"C2", X"DA", X"87", X"6A", X"3A", X"BB", --29D8
  X"61", X"D6", X"1E", X"38", X"05", X"D6", X"C2", X"DA", --29E0
  X"87", X"6A", X"CB", X"EE", X"C5", X"E5", X"3A", X"CC", --29E8
  X"61", X"D6", X"3E", X"38", X"0A", X"2A", X"AF", X"61", --29F0
  X"01", X"01", X"00", X"09", X"22", X"AF", X"61", X"E1", --29F8
  X"C1", X"3A", X"BA", X"61", X"D6", X"0A", X"38", X"04", --2A00
  X"D6", X"EA", X"38", X"31", X"3A", X"BB", X"61", X"D6", --2A08
  X"0A", X"38", X"04", X"D6", X"EA", X"38", X"26", X"CB", --2A10
  X"E6", X"3A", X"BA", X"61", X"D6", X"0A", X"30", X"06", --2A18
  X"CB", X"8E", X"CB", X"C6", X"18", X"04", X"CB", X"CE", --2A20
  X"CB", X"86", X"3A", X"BB", X"61", X"D6", X"0A", X"30", --2A28
  X"06", X"CB", X"96", X"CB", X"DE", X"18", X"50", X"CB", --2A30
  X"9E", X"CB", X"D6", X"18", X"4A", X"3A", X"BA", X"61", --2A38
  X"D6", X"0A", X"30", X"06", X"CB", X"8E", X"CB", X"86", --2A40
  X"18", X"18", X"D6", X"14", X"30", X"06", X"CB", X"C6", --2A48
  X"CB", X"8E", X"18", X"0E", X"D6", X"D6", X"30", X"06", --2A50
  X"CB", X"CE", X"CB", X"86", X"18", X"04", X"CB", X"8E", --2A58
  X"CB", X"86", X"3A", X"BB", X"61", X"D6", X"0A", X"30", --2A60
  X"06", X"CB", X"96", X"CB", X"9E", X"18", X"18", X"D6", --2A68
  X"14", X"30", X"06", X"CB", X"DE", X"CB", X"96", X"18", --2A70
  X"0E", X"D6", X"D6", X"30", X"06", X"CB", X"D6", X"CB", --2A78
  X"9E", X"18", X"04", X"CB", X"96", X"CB", X"9E", X"C9", --2A80
  X"21", X"5C", X"72", X"11", X"C0", X"61", X"3A", X"CC", --2A88
  X"61", X"96", X"38", X"19", X"23", X"96", X"30", X"16", --2A90
  X"23", X"3A", X"CB", X"61", X"96", X"38", X"10", X"23", --2A98
  X"96", X"30", X"0D", X"23", X"1A", X"E6", X"F0", X"4F", --2AA0
  X"7E", X"B1", X"12", X"18", X"09", X"23", X"23", X"23", --2AA8
  X"23", X"23", X"34", X"35", X"20", X"D8", X"C9", X"C9", --2AB0
  X"21", X"98", X"B7", X"11", X"00", X"40", X"ED", X"B0", --2AB8
  X"C9", X"01", X"00", X"03", X"21", X"30", X"75", X"11", --2AC0
  X"00", X"58", X"ED", X"B0", X"C9", X"F5", X"C5", X"3A", --2AC8
  X"78", X"5C", X"4F", X"3A", X"78", X"5C", X"91", X"28", --2AD0
  X"FA", X"C1", X"F1", X"C9", X"CD", X"CD", X"6A", X"CD", --2AD8
  X"E4", X"6A", X"18", X"0C", X"01", X"00", X"03", X"21", --2AE0
  X"31", X"78", X"11", X"00", X"58", X"ED", X"B0", X"C9", --2AE8
  X"CD", X"10", X"72", X"CD", X"CD", X"6A", X"CD", X"C1", --2AF0
  X"6A", X"CD", X"5A", X"71", X"C9", X"CD", X"CD", X"6A", --2AF8
  X"01", X"00", X"01", X"21", X"24", X"5E", X"11", X"C0", --2B00
  X"59", X"ED", X"B0", X"C9", X"01", X"C0", X"01", X"21", --2B08
  X"00", X"58", X"09", X"54", X"5D", X"21", X"30", X"75", --2B10
  X"09", X"01", X"00", X"01", X"ED", X"B0", X"C9", X"CD", --2B18
  X"FD", X"6A", X"CD", X"42", X"72", X"CD", X"CD", X"6A", --2B20
  X"CD", X"0C", X"6B", X"CD", X"5A", X"71", X"CD", X"F1", --2B28
  X"71", X"C9", X"01", X"28", X"00", X"21", X"F9", X"72", --2B30
  X"11", X"22", X"73", X"ED", X"B0", X"C9", X"21", X"DC", --2B38
  X"72", X"11", X"C0", X"61", X"1A", X"4F", X"CB", X"88", --2B40
  X"3A", X"CC", X"61", X"96", X"28", X"07", X"3C", X"3C", --2B48
  X"3D", X"28", X"02", X"18", X"08", X"CB", X"D9", X"CB", --2B50
  X"91", X"CB", X"C8", X"18", X"02", X"38", X"43", X"23", --2B58
  X"96", X"20", X"08", X"CB", X"99", X"CB", X"D1", X"CB", --2B60
  X"C8", X"18", X"02", X"30", X"36", X"23", X"3A", X"CB", --2B68
  X"61", X"96", X"20", X"08", X"CB", X"89", X"CB", X"C1", --2B70
  X"CB", X"C8", X"18", X"02", X"38", X"26", X"23", X"96", --2B78
  X"28", X"05", X"3D", X"28", X"02", X"18", X"08", X"CB", --2B80
  X"C9", X"CB", X"81", X"CB", X"C8", X"18", X"02", X"30", --2B88
  X"14", X"CB", X"48", X"28", X"03", X"79", X"12", X"C9", --2B90
  X"3A", X"C0", X"61", X"CB", X"FF", X"12", X"CD", X"41", --2B98
  X"6C", X"C9", X"23", X"23", X"23", X"23", X"34", X"35", --2BA0
  X"20", X"9E", X"C9", X"CB", X"90", X"3A", X"70", X"73", --2BA8
  X"21", X"76", X"72", X"3D", X"28", X"03", X"21", X"9F", --2BB0
  X"72", X"3A", X"C0", X"61", X"4F", X"CB", X"90", X"CB", --2BB8
  X"88", X"3A", X"CC", X"61", X"96", X"20", X"08", X"CB", --2BC0
  X"D1", X"CB", X"99", X"CB", X"C8", X"18", X"02", X"38", --2BC8
  X"5B", X"23", X"96", X"20", X"08", X"CB", X"D9", X"CB", --2BD0
  X"91", X"CB", X"C8", X"18", X"02", X"30", X"4E", X"23", --2BD8
  X"3A", X"CB", X"61", X"96", X"20", X"08", X"CB", X"C9", --2BE0
  X"CB", X"81", X"CB", X"C8", X"18", X"02", X"38", X"3E", --2BE8
  X"23", X"96", X"20", X"08", X"CB", X"C1", X"CB", X"89", --2BF0
  X"CB", X"C8", X"18", X"14", X"30", X"31", X"CB", X"48", --2BF8
  X"3A", X"73", X"73", X"23", X"96", X"20", X"09", X"21", --2C00
  X"C0", X"61", X"CB", X"FE", X"CD", X"36", X"6C", X"C9", --2C08
  X"11", X"C0", X"61", X"CB", X"48", X"28", X"07", X"79", --2C10
  X"CB", X"E7", X"CB", X"EF", X"12", X"C9", X"CB", X"D0", --2C18
  X"1A", X"E6", X"F0", X"4F", X"CD", X"A3", X"69", X"E6", --2C20
  X"0F", X"B1", X"12", X"C9", X"23", X"23", X"23", X"23", --2C28
  X"23", X"34", X"35", X"20", X"8A", X"C9", X"ED", X"4B", --2C30
  X"C5", X"61", X"CD", X"97", X"68", X"CD", X"DC", X"6A", --2C38
  X"C9", X"ED", X"4B", X"C5", X"61", X"CD", X"97", X"68", --2C40
  X"CD", X"1F", X"6B", X"C9", X"21", X"CB", X"61", X"3E", --2C48
  X"D8", X"77", X"21", X"CC", X"61", X"3E", X"A0", X"77", --2C50
  X"21", X"9D", X"6C", X"CD", X"83", X"6D", X"21", X"CB", --2C58
  X"61", X"3E", X"F0", X"77", X"21", X"9D", X"6C", X"CD", --2C60
  X"83", X"6D", X"3E", X"F8", X"21", X"CB", X"61", X"77", --2C68
  X"21", X"9D", X"6C", X"CD", X"83", X"6D", X"3E", X"AE", --2C70
  X"21", X"CC", X"61", X"77", X"21", X"CB", X"61", X"3E", --2C78
  X"D8", X"77", X"21", X"95", X"6C", X"CD", X"83", X"6D", --2C80
  X"21", X"CC", X"61", X"3E", X"A6", X"77", X"21", X"95", --2C88
  X"6C", X"CD", X"83", X"6D", X"C9", X"C0", X"00", X"80", --2C90
  X"00", X"C0", X"00", X"80", X"00", X"00", X"10", X"FF", --2C98
  X"10", X"10", X"FF", X"10", X"10", X"21", X"CB", X"61", --2CA0
  X"3E", X"E0", X"77", X"21", X"CC", X"61", X"3E", X"A0", --2CA8
  X"77", X"21", X"1E", X"6E", X"CD", X"83", X"6D", X"21", --2CB0
  X"CB", X"61", X"7E", X"C6", X"08", X"77", X"21", X"26", --2CB8
  X"6E", X"CD", X"83", X"6D", X"C9", X"21", X"CB", X"61", --2CC0
  X"3E", X"E8", X"77", X"21", X"CC", X"61", X"3E", X"A0", --2CC8
  X"77", X"21", X"2E", X"6E", X"CD", X"83", X"6D", X"21", --2CD0
  X"CC", X"61", X"7E", X"DE", X"08", X"77", X"21", X"36", --2CD8
  X"6E", X"CD", X"83", X"6D", X"C9", X"C9", X"3A", X"70", --2CE0
  X"73", X"11", X"A6", X"6D", X"3D", X"28", X"20", X"11", --2CE8
  X"DE", X"6D", X"3D", X"28", X"1A", X"CD", X"0F", X"6D", --2CF0
  X"11", X"16", X"6E", X"21", X"CC", X"61", X"3E", X"0F", --2CF8
  X"77", X"21", X"30", X"75", X"01", X"C0", X"02", X"09", --2D00
  X"22", X"A4", X"6D", X"0E", X"02", X"18", X"12", X"21", --2D08
  X"CC", X"61", X"3E", X"AF", X"77", X"21", X"30", X"75", --2D10
  X"01", X"40", X"00", X"09", X"22", X"A4", X"6D", X"0E", --2D18
  X"0E", X"C5", X"CD", X"31", X"6D", X"21", X"CC", X"61", --2D20
  X"7E", X"D6", X"08", X"77", X"C1", X"0D", X"20", X"F1", --2D28
  X"C9", X"01", X"04", X"00", X"21", X"CB", X"61", X"3E", --2D30
  X"00", X"77", X"C5", X"D5", X"CD", X"46", X"6D", X"D1", --2D38
  X"C1", X"13", X"0D", X"20", X"F5", X"C9", X"01", X"08", --2D40
  X"00", X"1A", X"C5", X"CB", X"7F", X"F5", X"28", X"09", --2D48
  X"CD", X"6E", X"6D", X"2A", X"A4", X"6D", X"3E", X"60", --2D50
  X"77", X"21", X"CB", X"61", X"7E", X"C6", X"08", X"77", --2D58
  X"2A", X"A4", X"6D", X"23", X"22", X"A4", X"6D", X"F1", --2D60
  X"17", X"C1", X"0D", X"20", X"DD", X"C9", X"CD", X"A3", --2D68
  X"69", X"E6", X"07", X"3C", X"21", X"46", X"6E", X"4F", --2D70
  X"0D", X"28", X"08", X"C5", X"01", X"08", X"00", X"09", --2D78
  X"C1", X"18", X"F5", X"22", X"C9", X"61", X"0E", X"08", --2D80
  X"2A", X"CB", X"61", X"E5", X"C5", X"CD", X"39", X"69", --2D88
  X"2A", X"C9", X"61", X"23", X"22", X"C9", X"61", X"21", --2D90
  X"CC", X"61", X"35", X"C1", X"0D", X"20", X"ED", X"E1", --2D98
  X"22", X"CB", X"61", X"C9", X"00", X"00", X"F0", X"00", --2DA0
  X"3F", X"80", X"F0", X"12", X"3F", X"00", X"C0", X"00", --2DA8
  X"1C", X"00", X"C0", X"00", X"0C", X"00", X"E0", X"00", --2DB0
  X"0E", X"03", X"C0", X"0C", X"0C", X"03", X"C0", X"3C", --2DB8
  X"00", X"0F", X"C0", X"7E", X"00", X"0F", X"E0", X"1C", --2DC0
  X"00", X"0F", X"E0", X"0C", X"00", X"0F", X"C0", X"0C", --2DC8
  X"00", X"0F", X"C0", X"0C", X"02", X"3F", X"C0", X"0C", --2DD0
  X"0F", X"FE", X"C0", X"0E", X"1D", X"DE", X"FF", X"86", --2DD8
  X"01", X"C0", X"C0", X"06", X"01", X"C0", X"E0", X"0E", --2DE0
  X"03", X"C0", X"C0", X"06", X"31", X"C3", X"C6", X"00", --2DE8
  X"30", X"03", X"C6", X"00", X"30", X"03", X"C6", X"60", --2DF0
  X"38", X"03", X"C6", X"7F", X"30", X"63", X"C6", X"7F", --2DF8
  X"30", X"63", X"C0", X"60", X"31", X"E0", X"C0", X"00", --2E00
  X"31", X"E0", X"80", X"00", X"F1", X"C0", X"00", X"01", --2E08
  X"F1", X"81", X"80", X"00", X"F0", X"03", X"E0", X"00", --2E10
  X"00", X"07", X"F0", X"00", X"00", X"17", X"80", X"FF", --2E18
  X"A0", X"84", X"FF", X"80", X"80", X"FF", X"01", X"FF", --2E20
  X"01", X"01", X"FF", X"21", X"05", X"FF", X"01", X"01", --2E28
  X"03", X"05", X"11", X"13", X"25", X"C9", X"92", X"A4", --2E30
  X"A8", X"90", X"A0", X"C0", X"80", X"00", X"18", X"7E", --2E38
  X"5E", X"FF", X"FF", X"7E", X"7E", X"18", X"10", X"38", --2E40
  X"54", X"38", X"54", X"BA", X"54", X"92", X"08", X"1C", --2E48
  X"2A", X"1C", X"2A", X"5D", X"2A", X"49", X"10", X"38", --2E50
  X"54", X"38", X"54", X"BA", X"54", X"10", X"08", X"1C", --2E58
  X"2A", X"1C", X"2A", X"5D", X"2A", X"08", X"00", X"10", --2E60
  X"38", X"54", X"38", X"54", X"10", X"10", X"10", X"38", --2E68
  X"54", X"38", X"54", X"10", X"10", X"00", X"00", X"04", --2E70
  X"0E", X"15", X"0E", X"15", X"04", X"04", X"04", X"0E", --2E78
  X"15", X"0E", X"15", X"04", X"04", X"00", X"3A", X"CB", --2E80
  X"61", X"D6", X"DC", X"D8", X"3A", X"CC", X"61", X"D6", --2E88
  X"92", X"D8", X"21", X"AB", X"61", X"CB", X"FE", X"21", --2E90
  X"C0", X"61", X"CB", X"FE", X"ED", X"4B", X"C5", X"61", --2E98
  X"CD", X"97", X"68", X"2A", X"CB", X"61", X"E5", X"2A", --2EA0
  X"C9", X"61", X"E5", X"CD", X"A5", X"6C", X"CD", X"C5", --2EA8
  X"6C", X"21", X"B5", X"61", X"34", X"2A", X"AF", X"61", --2EB0
  X"01", X"F4", X"01", X"09", X"22", X"AF", X"61", X"21", --2EB8
  X"F4", X"01", X"11", X"06", X"00", X"CD", X"32", X"72", --2EC0
  X"3A", X"B3", X"61", X"21", X"CB", X"61", X"77", X"D6", --2EC8
  X"08", X"21", X"B3", X"61", X"77", X"D6", X"D5", X"30", --2ED0
  X"09", X"3E", X"F7", X"77", X"21", X"B4", X"61", X"3E", --2ED8
  X"A8", X"77", X"3A", X"B3", X"61", X"21", X"CB", X"61", --2EE0
  X"77", X"3A", X"B4", X"61", X"21", X"CC", X"61", X"77", --2EE8
  X"01", X"D8", X"74", X"CD", X"97", X"68", X"CD", X"3A", --2EF0
  X"64", X"21", X"F4", X"01", X"11", X"03", X"00", X"CD", --2EF8
  X"32", X"72", X"CD", X"C5", X"6C", X"CD", X"A5", X"6C", --2F00
  X"E1", X"22", X"C9", X"61", X"E1", X"22", X"CB", X"61", --2F08
  X"C9", X"3A", X"73", X"73", X"3C", X"3D", X"C0", X"3A", --2F10
  X"CB", X"61", X"21", X"6F", X"73", X"96", X"C6", X"08", --2F18
  X"D6", X"10", X"D0", X"3A", X"CC", X"61", X"21", X"6E", --2F20
  X"73", X"96", X"C6", X"08", X"D6", X"10", X"D0", X"21", --2F28
  X"C0", X"61", X"CB", X"FE", X"CD", X"36", X"6C", X"C9", --2F30
  X"01", X"16", X"48", X"7F", X"20", X"42", X"55", X"4C", --2F38
  X"4C", X"41", X"52", X"01", X"39", X"48", X"31", X"39", --2F40
  X"38", X"34", X"01", X"00", X"48", X"4E", X"20", X"55", --2F48
  X"50", X"01", X"20", X"48", X"4D", X"20", X"44", X"4F", --2F50
  X"57", X"4E", X"01", X"40", X"48", X"5A", X"20", X"4C", --2F58
  X"45", X"46", X"54", X"01", X"60", X"48", X"58", X"20", --2F60
  X"52", X"49", X"47", X"48", X"54", X"01", X"8A", X"48", --2F68
  X"53", X"43", X"4F", X"52", X"45", X"01", X"AA", X"48", --2F70
  X"48", X"49", X"47", X"48", X"01", X"E9", X"48", X"53", --2F78
  X"50", X"41", X"43", X"45", X"20", X"54", X"4F", X"20", --2F80
  X"53", X"54", X"41", X"52", X"54", X"00", X"18", X"03", --2F88
  X"CD", X"47", X"70", X"21", X"D2", X"61", X"CB", X"E6", --2F90
  X"CB", X"AE", X"3E", X"7F", X"DB", X"FE", X"CB", X"57", --2F98
  X"20", X"15", X"3A", X"D4", X"61", X"D6", X"06", X"38", --2FA0
  X"2A", X"21", X"CD", X"61", X"CB", X"C6", X"CB", X"8E", --2FA8
  X"21", X"D4", X"61", X"35", X"35", X"18", X"1C", X"3E", --2FB0
  X"7F", X"DB", X"FE", X"CB", X"5F", X"00", X"20", X"13", --2FB8
  X"3A", X"D4", X"61", X"D6", X"AE", X"30", X"0C", X"21", --2FC0
  X"CD", X"61", X"CB", X"C6", X"CB", X"8E", X"21", X"D4", --2FC8
  X"61", X"34", X"34", X"3E", X"FE", X"00", X"DB", X"FE", --2FD0
  X"CB", X"57", X"00", X"20", X"1D", X"3A", X"D5", X"61", --2FD8
  X"D6", X"ED", X"D2", X"1E", X"70", X"21", X"D2", X"61", --2FE0
  X"CB", X"B6", X"CB", X"FE", X"21", X"CD", X"61", X"CB", --2FE8
  X"C6", X"CB", X"8E", X"21", X"D5", X"61", X"34", X"34", --2FF0
  X"18", X"24", X"3E", X"FE", X"DB", X"FE", X"CB", X"4F", --2FF8
  X"00", X"00", X"20", X"1A", X"3A", X"D5", X"61", X"D6", --3000
  X"02", X"38", X"13", X"21", X"D2", X"61", X"CB", X"F6", --3008
  X"CB", X"BE", X"21", X"CD", X"61", X"CB", X"C6", X"CB", --3010
  X"8E", X"21", X"D5", X"61", X"35", X"35", X"3A", X"70", --3018
  X"73", X"D6", X"04", X"30", X"03", X"CD", X"CD", X"6A", --3020
  X"21", X"CD", X"61", X"CB", X"46", X"20", X"11", X"CB", --3028
  X"4E", X"20", X"0C", X"CB", X"CE", X"21", X"D2", X"61", --3030
  X"CB", X"A6", X"CB", X"AE", X"CD", X"8C", X"70", X"C9", --3038
  X"CB", X"86", X"CD", X"7E", X"70", X"18", X"F8", X"01", --3040
  X"88", X"74", X"ED", X"43", X"D2", X"61", X"ED", X"43", --3048
  X"CE", X"61", X"01", X"10", X"40", X"ED", X"43", X"D4", --3050
  X"61", X"ED", X"43", X"D0", X"61", X"CD", X"AF", X"70", --3058
  X"C9", X"2A", X"D2", X"61", X"ED", X"4B", X"CE", X"61", --3060
  X"22", X"CE", X"61", X"ED", X"43", X"D2", X"61", X"2A", --3068
  X"D4", X"61", X"ED", X"4B", X"D0", X"61", X"22", X"D0", --3070
  X"61", X"ED", X"43", X"D4", X"61", X"C9", X"21", X"78", --3078
  X"5C", X"CB", X"5E", X"20", X"07", X"21", X"D2", X"61", --3080
  X"3E", X"30", X"AE", X"77", X"CD", X"AF", X"70", X"CD", --3088
  X"61", X"70", X"CD", X"AF", X"70", X"CD", X"61", X"70", --3090
  X"CD", X"5A", X"71", X"ED", X"4B", X"D2", X"61", X"ED", --3098
  X"43", X"CE", X"61", X"ED", X"4B", X"D4", X"61", X"ED", --30A0
  X"43", X"D0", X"61", X"CD", X"C6", X"71", X"C9", X"2A", --30A8
  X"D2", X"61", X"E5", X"2A", X"D4", X"61", X"E5", X"0E", --30B0
  X"05", X"C5", X"CD", X"D3", X"70", X"21", X"D2", X"61", --30B8
  X"34", X"34", X"21", X"D4", X"61", X"35", X"C1", X"0D", --30C0
  X"20", X"EF", X"E1", X"22", X"D4", X"61", X"E1", X"22", --30C8
  X"D2", X"61", X"C9", X"3A", X"D4", X"61", X"C6", X"08", --30D0
  X"F5", X"0F", X"0F", X"0F", X"E6", X"1F", X"47", X"3E", --30D8
  X"18", X"98", X"47", X"3A", X"D5", X"61", X"0F", X"0F", --30E0
  X"0F", X"E6", X"1F", X"4F", X"F1", X"E6", X"07", X"5F", --30E8
  X"3E", X"07", X"9B", X"CD", X"47", X"71", X"3A", X"D5", --30F0
  X"61", X"E6", X"07", X"4F", X"0C", X"0D", X"28", X"3A", --30F8
  X"3E", X"FF", X"C5", X"1F", X"CB", X"BF", X"0D", X"20", --3100
  X"FA", X"57", X"ED", X"4B", X"D2", X"61", X"0A", X"C1", --3108
  X"C5", X"0F", X"0D", X"20", X"FC", X"5F", X"A2", X"AE", --3110
  X"77", X"23", X"3E", X"FF", X"AA", X"57", X"7B", X"A2", --3118
  X"AE", X"77", X"ED", X"4B", X"D2", X"61", X"03", X"0A", --3120
  X"C1", X"0F", X"0D", X"20", X"FC", X"5F", X"3E", X"FF", --3128
  X"AA", X"A3", X"AE", X"77", X"7B", X"A2", X"23", X"AE", --3130
  X"77", X"C9", X"ED", X"4B", X"D2", X"61", X"0A", X"AE", --3138
  X"77", X"03", X"23", X"0A", X"AE", X"77", X"C9", X"F5", --3140
  X"78", X"E6", X"18", X"F6", X"40", X"67", X"F1", X"84", --3148
  X"67", X"78", X"E6", X"07", X"0F", X"0F", X"0F", X"81", --3150
  X"6F", X"C9", X"3A", X"D5", X"61", X"1F", X"1F", X"1F", --3158
  X"E6", X"1F", X"4F", X"AF", X"47", X"6F", X"67", X"3A", --3160
  X"D4", X"61", X"5F", X"3E", X"BF", X"93", X"E6", X"F8", --3168
  X"6F", X"CB", X"15", X"CB", X"14", X"AF", X"CB", X"15", --3170
  X"CB", X"14", X"09", X"01", X"00", X"58", X"09", X"E5", --3178
  X"ED", X"5B", X"B8", X"61", X"21", X"30", X"75", X"01", --3180
  X"00", X"58", X"ED", X"42", X"19", X"01", X"03", X"00", --3188
  X"ED", X"B0", X"3A", X"D4", X"61", X"D6", X"08", X"38", --3190
  X"10", X"01", X"1D", X"00", X"09", X"E5", X"6B", X"62", --3198
  X"09", X"5D", X"54", X"E1", X"01", X"03", X"00", X"ED", --31A0
  X"B0", X"E1", X"22", X"B8", X"61", X"3E", X"60", X"77", --31A8
  X"23", X"77", X"23", X"77", X"3A", X"D4", X"61", X"D6", --31B0
  X"08", X"D8", X"3E", X"60", X"01", X"1E", X"00", X"09", --31B8
  X"77", X"23", X"77", X"23", X"77", X"C9", X"3A", X"78", --31C0
  X"5C", X"CB", X"5F", X"21", X"CD", X"61", X"28", X"12", --31C8
  X"CB", X"7E", X"C0", X"CB", X"FE", X"11", X"01", X"00", --31D0
  X"21", X"C2", X"01", X"CD", X"B5", X"03", X"CD", X"3A", --31D8
  X"64", X"C9", X"CB", X"7E", X"C8", X"CB", X"BE", X"11", --31E0
  X"01", X"00", X"21", X"90", X"01", X"CD", X"B5", X"03", --31E8
  X"C9", X"21", X"FA", X"00", X"CD", X"2F", X"72", X"21", --31F0
  X"C2", X"01", X"CD", X"2F", X"72", X"21", X"90", X"01", --31F8
  X"CD", X"2F", X"72", X"21", X"5E", X"01", X"CD", X"2F", --3200
  X"72", X"21", X"2C", X"01", X"CD", X"2F", X"72", X"C9", --3208
  X"21", X"58", X"02", X"11", X"02", X"00", X"CD", X"32", --3210
  X"72", X"11", X"0A", X"00", X"21", X"2C", X"01", X"0E", --3218
  X"50", X"E5", X"D5", X"C5", X"CD", X"B5", X"03", X"C1", --3220
  X"D1", X"E1", X"23", X"0D", X"20", X"F3", X"C9", X"11", --3228
  X"03", X"00", X"E5", X"D5", X"CD", X"B5", X"03", X"D1", --3230
  X"E1", X"01", X"08", X"00", X"AF", X"ED", X"42", X"30", --3238
  X"F1", X"C9", X"0E", X"C8", X"C5", X"CD", X"A3", X"69", --3240
  X"6F", X"E6", X"03", X"67", X"3E", X"01", X"5F", X"3E", --3248
  X"00", X"57", X"CD", X"B5", X"03", X"C1", X"0D", X"C5", --3250
  X"20", X"EB", X"C1", X"C9", X"34", X"06", X"2C", X"0D", --3258
  X"06", X"18", X"1C", X"2D", X"0A", X"04", X"20", X"12", --3260
  X"14", X"18", X"02", X"A0", X"10", X"EC", X"10", X"06", --3268
  X"98", X"20", X"D2", X"14", X"09", X"00", X"40", X"64", --3270
  X"01", X"0A", X"01", X"A4", X"0A", X"01", X"1B", X"01", --3278
  X"44", X"48", X"5C", X"10", X"02", X"74", X"10", X"50", --3280
  X"20", X"02", X"A4", X"0A", X"8C", X"30", X"03", X"84", --3288
  X"20", X"9C", X"10", X"03", X"44", X"10", X"9C", X"60", --3290
  X"04", X"44", X"40", X"DC", X"20", X"04", X"00", X"5C", --3298
  X"58", X"01", X"0A", X"01", X"AE", X"08", X"0A", X"38", --32A0
  X"01", X"74", X"20", X"24", X"10", X"02", X"64", X"20", --32A8
  X"44", X"10", X"03", X"6C", X"10", X"44", X"40", X"03", --32B0
  X"94", X"20", X"64", X"10", X"04", X"44", X"18", X"7C", --32B8
  X"20", X"05", X"44", X"58", X"8C", X"10", X"05", X"94", --32C0
  X"20", X"B4", X"18", X"06", X"4C", X"18", X"B4", X"10", --32C8
  X"07", X"5C", X"20", X"C4", X"10", X"07", X"6C", X"18", --32D0
  X"EC", X"0E", X"08", X"00", X"14", X"30", X"01", X"13", --32D8
  X"34", X"06", X"14", X"18", X"34", X"06", X"3C", X"22", --32E0
  X"29", X"0B", X"5C", X"08", X"24", X"06", X"5C", X"68", --32E8
  X"29", X"13", X"BC", X"08", X"3C", X"05", X"BC", X"41", --32F0
  X"00", X"DA", X"14", X"00", X"00", X"DC", X"0A", X"00", --32F8
  X"00", X"DA", X"10", X"00", X"00", X"D2", X"10", X"00", --3300
  X"00", X"DE", X"19", X"00", X"00", X"D8", X"18", X"00", --3308
  X"00", X"D2", X"0E", X"00", X"00", X"D2", X"1E", X"00", --3310
  X"00", X"D7", X"14", X"00", X"00", X"D8", X"20", X"00", --3318
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3320
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3328
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3330
  X"00", X"00", X"00", X"00", X"10", X"D0", X"05", X"E3", --3338
  X"1E", X"D8", X"06", X"D4", X"1B", X"D0", X"08", X"CF", --3340
  X"0D", X"D0", X"05", X"D0", X"1F", X"D0", X"05", X"D4", --3348
  X"13", X"D0", X"05", X"D8", X"23", X"D8", X"08", X"00", --3350
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3358
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3360
  X"00", X"00", X"00", X"00", X"00", X"00", X"47", X"82", --3368
  X"01", X"3E", X"00", X"FF", X"00", X"00", X"00", X"00", --3370
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3378
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3380
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3388
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3390
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3398
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --33A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --33A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --33B0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --33B8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --33C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --33C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --33D0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --33D8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --33E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --33E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --33F0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --33F8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3400
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3408
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3410
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3418
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3420
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3428
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3430
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3438
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3440
  X"00", X"00", X"08", X"00", X"3F", X"FC", X"0F", X"F3", --3448
  X"79", X"E0", X"00", X"E1", X"00", X"00", X"00", X"00", --3450
  X"08", X"00", X"3F", X"FC", X"0F", X"F3", X"18", X"30", --3458
  X"20", X"08", X"00", X"00", X"00", X"00", X"00", X"00", --3460
  X"08", X"03", X"3F", X"FC", X"0F", X"E0", X"04", X"60", --3468
  X"02", X"80", X"00", X"00", X"00", X"00", X"0C", X"00", --3470
  X"3F", X"FC", X"07", X"F2", X"06", X"31", X"04", X"10", --3478
  X"0C", X"30", X"00", X"00", X"00", X"00", X"00", X"00", --3480
  X"00", X"00", X"00", X"10", X"3F", X"FC", X"CF", X"F0", --3488
  X"07", X"9E", X"00", X"00", X"00", X"00", X"00", X"00", --3490
  X"00", X"10", X"3F", X"FC", X"CF", X"F0", X"0C", X"30", --3498
  X"10", X"08", X"00", X"00", X"00", X"00", X"00", X"00", --34A0
  X"C0", X"10", X"3F", X"FC", X"0F", X"F0", X"0C", X"20", --34A8
  X"02", X"40", X"3A", X"EF", X"7E", X"47", X"01", X"80", --34B0
  X"3E", X"4C", X"D8", X"49", X"4A", X"D8", X"56", X"47", --34B8
  X"D8", X"61", X"44", X"D8", X"69", X"46", X"D8", X"4B", --34C0
  X"51", X"D8", X"55", X"52", X"D8", X"5D", X"53", X"D8", --34C8
  X"3E", X"FF", X"FF", X"7F", X"22", X"22", X"1F", X"00", --34D0
  X"7C", X"FF", X"FF", X"FE", X"44", X"44", X"23", X"10", --34D8
  X"FB", X"11", X"E0", X"00", X"78", X"7F", X"0A", X"01", --34E0
  X"03", X"0A", X"0A", X"03", X"00", X"D8", X"FF", X"91", --34E8
  X"52", X"D8", X"FF", X"91", X"52", X"E2", X"88", X"FF", --34F0
  X"4E", X"46", X"98", X"FF", X"4E", X"46", X"3C", X"00", --34F8
  X"F3", X"AF", X"11", X"FF", X"FF", X"C3", X"CB", X"11", --3500
  X"2A", X"5D", X"5C", X"22", X"5F", X"5C", X"18", X"43", --3508
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3510
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3518
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3520
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3528
  X"75", X"75", X"65", X"65", X"65", X"65", X"65", X"65", --3530
  X"65", X"65", X"65", X"65", X"65", X"65", X"65", X"65", --3538
  X"65", X"65", X"65", X"65", X"65", X"65", X"7D", X"7D", --3540
  X"78", X"78", X"78", X"78", X"78", X"78", X"7D", X"7D", --3548
  X"75", X"75", X"65", X"65", X"65", X"65", X"65", X"65", --3550
  X"65", X"65", X"65", X"65", X"65", X"65", X"65", X"65", --3558
  X"65", X"65", X"65", X"65", X"65", X"65", X"65", X"7D", --3560
  X"7D", X"7D", X"7D", X"7D", X"7D", X"7D", X"7D", X"65", --3568
  X"60", X"60", X"60", X"60", X"67", X"67", X"67", X"67", --3570
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3578
  X"67", X"67", X"60", X"60", X"60", X"60", X"60", X"60", --3580
  X"60", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3588
  X"60", X"60", X"60", X"60", X"67", X"67", X"67", X"67", --3590
  X"67", X"67", X"67", X"60", X"67", X"67", X"60", X"67", --3598
  X"67", X"67", X"60", X"60", X"60", X"60", X"60", X"60", --35A0
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --35A8
  X"60", X"60", X"67", X"67", X"67", X"67", X"67", X"67", --35B0
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --35B8
  X"67", X"67", X"67", X"60", X"60", X"60", X"67", X"67", --35C0
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --35C8
  X"60", X"60", X"67", X"67", X"67", X"67", X"67", X"67", --35D0
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --35D8
  X"67", X"67", X"67", X"67", X"60", X"60", X"67", X"67", --35E0
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --35E8
  X"60", X"60", X"60", X"67", X"67", X"67", X"67", X"67", --35F0
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --35F8
  X"67", X"67", X"67", X"67", X"60", X"60", X"60", X"67", --3600
  X"67", X"67", X"67", X"67", X"67", X"67", X"60", X"60", --3608
  X"60", X"60", X"67", X"67", X"67", X"67", X"67", X"67", --3610
  X"67", X"67", X"67", X"67", X"60", X"60", X"67", X"67", --3618
  X"67", X"67", X"67", X"67", X"60", X"60", X"67", X"67", --3620
  X"67", X"67", X"67", X"67", X"67", X"67", X"60", X"60", --3628
  X"60", X"60", X"67", X"67", X"67", X"67", X"67", X"67", --3630
  X"67", X"67", X"60", X"60", X"60", X"60", X"67", X"67", --3638
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3640
  X"67", X"67", X"67", X"67", X"60", X"60", X"60", X"60", --3648
  X"60", X"60", X"67", X"67", X"67", X"67", X"67", X"67", --3650
  X"67", X"60", X"60", X"60", X"60", X"60", X"60", X"67", --3658
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3660
  X"67", X"67", X"67", X"67", X"60", X"60", X"60", X"60", --3668
  X"60", X"60", X"60", X"67", X"67", X"67", X"67", X"67", --3670
  X"67", X"67", X"67", X"60", X"60", X"60", X"67", X"67", --3678
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3680
  X"67", X"67", X"67", X"67", X"60", X"60", X"60", X"60", --3688
  X"60", X"60", X"60", X"67", X"67", X"67", X"67", X"67", --3690
  X"67", X"67", X"67", X"67", X"60", X"60", X"67", X"67", --3698
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --36A0
  X"67", X"67", X"67", X"67", X"60", X"60", X"60", X"60", --36A8
  X"60", X"60", X"67", X"67", X"67", X"67", X"67", X"67", --36B0
  X"67", X"67", X"67", X"67", X"60", X"60", X"67", X"67", --36B8
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --36C0
  X"67", X"67", X"67", X"67", X"60", X"60", X"60", X"60", --36C8
  X"60", X"60", X"67", X"67", X"67", X"67", X"67", X"67", --36D0
  X"67", X"67", X"67", X"67", X"60", X"60", X"67", X"67", --36D8
  X"67", X"67", X"67", X"67", X"67", X"67", X"60", X"67", --36E0
  X"67", X"67", X"60", X"60", X"60", X"60", X"60", X"60", --36E8
  X"60", X"60", X"67", X"67", X"67", X"67", X"67", X"67", --36F0
  X"67", X"67", X"67", X"67", X"60", X"60", X"67", X"67", --36F8
  X"67", X"67", X"67", X"67", X"60", X"60", X"60", X"60", --3700
  X"60", X"60", X"60", X"60", X"60", X"60", X"60", X"67", --3708
  X"60", X"60", X"67", X"67", X"67", X"67", X"67", X"67", --3710
  X"67", X"67", X"67", X"67", X"60", X"60", X"60", X"67", --3718
  X"67", X"67", X"67", X"60", X"60", X"60", X"67", X"60", --3720
  X"60", X"60", X"67", X"60", X"60", X"60", X"60", X"67", --3728
  X"61", X"61", X"61", X"67", X"67", X"67", X"67", X"67", --3730
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3738
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3740
  X"61", X"61", X"61", X"61", X"61", X"61", X"61", X"61", --3748
  X"61", X"61", X"61", X"61", X"61", X"61", X"67", X"67", --3750
  X"61", X"61", X"61", X"61", X"61", X"67", X"67", X"67", --3758
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3760
  X"61", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3768
  X"61", X"61", X"61", X"67", X"67", X"67", X"67", X"67", --3770
  X"67", X"67", X"67", X"67", X"61", X"67", X"67", X"67", --3778
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3780
  X"61", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3788
  X"61", X"61", X"61", X"67", X"67", X"67", X"67", X"67", --3790
  X"67", X"67", X"67", X"67", X"61", X"61", X"61", X"61", --3798
  X"61", X"61", X"61", X"61", X"61", X"61", X"61", X"61", --37A0
  X"61", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --37A8
  X"61", X"61", X"61", X"67", X"67", X"67", X"67", X"67", --37B0
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --37B8
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --37C0
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --37C8
  X"61", X"61", X"61", X"67", X"67", X"67", X"67", X"67", --37D0
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --37D8
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --37E0
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --37E8
  X"60", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --37F0
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --37F8
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3800
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3808
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3810
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3818
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3820
  X"67", X"67", X"67", X"67", X"67", X"67", X"67", X"67", --3828
  X"67", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3830
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3838
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3840
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3848
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3850
  X"00", X"52", X"00", X"00", X"00", X"00", X"00", X"00", --3858
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3860
  X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3868
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3870
  X"00", X"52", X"52", X"00", X"00", X"00", X"00", X"00", --3878
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", --3880
  X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3888
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3890
  X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", --3898
  X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", --38A0
  X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", --38A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --38B0
  X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"12", --38B8
  X"12", X"12", X"12", X"00", X"00", X"00", X"52", X"52", --38C0
  X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", --38C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --38D0
  X"52", X"52", X"52", X"52", X"52", X"52", X"12", X"12", --38D8
  X"12", X"12", X"12", X"12", X"52", X"52", X"52", X"52", --38E0
  X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", --38E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --38F0
  X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"12", --38F8
  X"12", X"12", X"12", X"52", X"52", X"52", X"52", X"52", --3900
  X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", --3908
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3910
  X"00", X"52", X"52", X"52", X"76", X"76", X"52", X"52", --3918
  X"12", X"12", X"52", X"52", X"76", X"76", X"52", X"52", --3920
  X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3928
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3930
  X"00", X"52", X"52", X"76", X"00", X"76", X"76", X"52", --3938
  X"12", X"12", X"52", X"76", X"00", X"76", X"76", X"52", --3940
  X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3948
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3950
  X"00", X"52", X"52", X"52", X"76", X"76", X"52", X"52", --3958
  X"12", X"12", X"52", X"52", X"76", X"76", X"52", X"52", --3960
  X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3968
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3970
  X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", --3978
  X"12", X"12", X"52", X"52", X"52", X"52", X"52", X"52", --3980
  X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3988
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3990
  X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", --3998
  X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", --39A0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --39A8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --39B0
  X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"00", --39B8
  X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", --39C0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --39C8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --39D0
  X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"00", --39D8
  X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", --39E0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --39E8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --39F0
  X"00", X"00", X"00", X"52", X"52", X"52", X"12", X"7F", --39F8
  X"12", X"12", X"7F", X"12", X"52", X"52", X"52", X"00", --3A00
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3A08
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3A10
  X"00", X"00", X"00", X"00", X"52", X"52", X"12", X"7F", --3A18
  X"12", X"12", X"7F", X"12", X"52", X"52", X"00", X"00", --3A20
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3A28
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3A30
  X"00", X"00", X"00", X"00", X"00", X"12", X"12", X"7F", --3A38
  X"12", X"12", X"7F", X"12", X"12", X"00", X"00", X"00", --3A40
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3A48
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3A50
  X"00", X"00", X"00", X"00", X"00", X"12", X"12", X"12", --3A58
  X"12", X"12", X"12", X"12", X"12", X"00", X"00", X"00", --3A60
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3A68
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3A70
  X"00", X"00", X"00", X"00", X"00", X"00", X"12", X"12", --3A78
  X"12", X"12", X"12", X"12", X"00", X"00", X"00", X"00", --3A80
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3A88
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3A90
  X"00", X"00", X"00", X"00", X"00", X"00", X"12", X"7F", --3A98
  X"12", X"12", X"7F", X"12", X"00", X"00", X"00", X"00", --3AA0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3AA8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3AB0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"7F", --3AB8
  X"12", X"12", X"7F", X"00", X"00", X"00", X"00", X"00", --3AC0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3AC8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3AD0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", --3AD8
  X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", --3AE0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3AE8
  X"00", X"07", X"07", X"07", X"07", X"07", X"07", X"07", --3AF0
  X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", --3AF8
  X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", --3B00
  X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", --3B08
  X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", --3B10
  X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", --3B18
  X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", --3B20
  X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", --3B28
  X"07", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3B30
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3B38
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3B40
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3B48
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3B50
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3B58
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3B60
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3B68
  X"18", X"2F", X"C3", X"88", X"7B", X"00", X"00", X"00", --3B70
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3B78
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3B80
  X"21", X"02", X"00", X"22", X"86", X"7B", X"3E", X"1E", --3B88
  X"21", X"84", X"7B", X"77", X"3E", X"00", X"21", X"77", --3B90
  X"7B", X"77", X"3E", X"01", X"21", X"75", X"7B", X"77", --3B98
  X"C9", X"3A", X"77", X"7B", X"3C", X"3D", X"28", X"15", --3BA0
  X"3D", X"3D", X"20", X"11", X"CD", X"49", X"7F", X"CD", --3BA8
  X"91", X"7C", X"21", X"77", X"7B", X"35", X"35", X"21", --3BB0
  X"72", X"73", X"CB", X"CE", X"C9", X"3A", X"77", X"7B", --3BB8
  X"3C", X"3D", X"C2", X"6F", X"7C", X"21", X"84", X"7B", --3BC0
  X"35", X"28", X"12", X"21", X"73", X"73", X"3E", X"FF", --3BC8
  X"77", X"3A", X"84", X"7B", X"D6", X"05", X"30", X"04", --3BD0
  X"3A", X"75", X"7B", X"77", X"C9", X"3E", X"1E", X"77", --3BD8
  X"3A", X"70", X"73", X"21", X"89", X"7E", X"3D", X"28", --3BE0
  X"33", X"21", X"C9", X"7E", X"3D", X"28", X"2D", X"3A", --3BE8
  X"75", X"7B", X"3D", X"20", X"27", X"3A", X"71", X"73", --3BF0
  X"CB", X"5F", X"20", X"20", X"11", X"6F", X"73", X"3E", --3BF8
  X"01", X"12", X"11", X"6E", X"73", X"3E", X"07", X"12", --3C00
  X"11", X"79", X"7B", X"3E", X"02", X"12", X"11", X"76", --3C08
  X"7B", X"3E", X"E0", X"12", X"11", X"75", X"7B", X"3E", --3C10
  X"08", X"12", X"18", X"3B", X"3E", X"00", X"47", X"3A", --3C18
  X"75", X"7B", X"3D", X"CB", X"07", X"4F", X"3A", X"71", --3C20
  X"73", X"CB", X"4F", X"20", X"01", X"0C", X"79", X"CB", --3C28
  X"07", X"CB", X"07", X"CB", X"07", X"4F", X"09", X"7E", --3C30
  X"23", X"11", X"6F", X"73", X"12", X"7E", X"23", X"11", --3C38
  X"6E", X"73", X"3D", X"12", X"7E", X"23", X"11", X"79", --3C40
  X"7B", X"12", X"7E", X"23", X"11", X"76", X"7B", X"D6", --3C48
  X"10", X"12", X"7E", X"11", X"75", X"7B", X"12", X"CD", --3C50
  X"91", X"7C", X"3A", X"76", X"7B", X"21", X"77", X"7B", --3C58
  X"77", X"21", X"82", X"7B", X"3A", X"76", X"7B", X"CB", --3C60
  X"0F", X"CB", X"0F", X"CB", X"0F", X"77", X"C9", X"21", --3C68
  X"73", X"73", X"3E", X"00", X"77", X"21", X"6F", X"73", --3C70
  X"3A", X"79", X"7B", X"CB", X"4F", X"20", X"04", X"35", --3C78
  X"35", X"18", X"02", X"34", X"34", X"CD", X"C1", X"7C", --3C80
  X"CD", X"C9", X"7D", X"21", X"77", X"7B", X"35", X"35", --3C88
  X"C9", X"CD", X"1E", X"7E", X"2A", X"80", X"7B", X"22", --3C90
  X"7C", X"7B", X"2A", X"6E", X"73", X"22", X"7E", X"7B", --3C98
  X"CD", X"1E", X"7D", X"C9", X"2A", X"80", X"7B", X"ED", --3CA0
  X"4B", X"7C", X"7B", X"22", X"7C", X"7B", X"ED", X"43", --3CA8
  X"80", X"7B", X"2A", X"6E", X"73", X"ED", X"4B", X"7E", --3CB0
  X"7B", X"22", X"7E", X"7B", X"ED", X"43", X"6E", X"73", --3CB8
  X"C9", X"CD", X"1E", X"7E", X"CD", X"D8", X"7C", X"ED", --3CC0
  X"4B", X"80", X"7B", X"ED", X"43", X"7C", X"7B", X"ED", --3CC8
  X"4B", X"6E", X"73", X"ED", X"43", X"7E", X"7B", X"C9", --3CD0
  X"2A", X"80", X"7B", X"E5", X"2A", X"6E", X"73", X"E5", --3CD8
  X"2A", X"7C", X"7B", X"E5", X"2A", X"7E", X"7B", X"E5", --3CE0
  X"0E", X"08", X"C5", X"CD", X"42", X"7D", X"21", X"80", --3CE8
  X"7B", X"34", X"34", X"21", X"6E", X"73", X"35", X"CD", --3CF0
  X"A4", X"7C", X"CD", X"42", X"7D", X"21", X"80", X"7B", --3CF8
  X"34", X"34", X"21", X"6E", X"73", X"35", X"CD", X"A4", --3D00
  X"7C", X"C1", X"0D", X"20", X"DD", X"E1", X"22", X"7E", --3D08
  X"7B", X"E1", X"22", X"7C", X"7B", X"E1", X"22", X"6E", --3D10
  X"73", X"E1", X"22", X"80", X"7B", X"C9", X"2A", X"80", --3D18
  X"7B", X"E5", X"2A", X"6E", X"73", X"E5", X"0E", X"08", --3D20
  X"C5", X"CD", X"42", X"7D", X"21", X"80", X"7B", X"34", --3D28
  X"34", X"21", X"6E", X"73", X"35", X"C1", X"0D", X"20", --3D30
  X"EF", X"E1", X"22", X"6E", X"73", X"E1", X"22", X"80", --3D38
  X"7B", X"C9", X"3A", X"6E", X"73", X"C6", X"08", X"F5", --3D40
  X"0F", X"0F", X"0F", X"E6", X"1F", X"47", X"3E", X"18", --3D48
  X"98", X"47", X"3A", X"6F", X"73", X"0F", X"0F", X"0F", --3D50
  X"E6", X"1F", X"4F", X"F1", X"E6", X"07", X"5F", X"3E", --3D58
  X"07", X"9B", X"CD", X"B6", X"7D", X"3A", X"6F", X"73", --3D60
  X"E6", X"07", X"4F", X"0C", X"0D", X"28", X"3A", X"3E", --3D68
  X"FF", X"C5", X"1F", X"CB", X"BF", X"0D", X"20", X"FA", --3D70
  X"57", X"ED", X"4B", X"80", X"7B", X"0A", X"C1", X"C5", --3D78
  X"0F", X"0D", X"20", X"FC", X"5F", X"A2", X"AE", X"77", --3D80
  X"23", X"3E", X"FF", X"AA", X"57", X"7B", X"A2", X"AE", --3D88
  X"77", X"ED", X"4B", X"80", X"7B", X"03", X"0A", X"C1", --3D90
  X"0F", X"0D", X"20", X"FC", X"5F", X"3E", X"FF", X"AA", --3D98
  X"A3", X"AE", X"77", X"7B", X"A2", X"23", X"AE", X"77", --3DA0
  X"C9", X"ED", X"4B", X"80", X"7B", X"0A", X"AE", X"77", --3DA8
  X"03", X"23", X"0A", X"AE", X"77", X"C9", X"F5", X"78", --3DB0
  X"E6", X"18", X"F6", X"40", X"67", X"F1", X"84", X"67", --3DB8
  X"78", X"E6", X"07", X"0F", X"0F", X"0F", X"81", X"6F", --3DC0
  X"C9", X"CD", X"49", X"7F", X"3A", X"6F", X"73", X"1F", --3DC8
  X"1F", X"1F", X"E6", X"1F", X"4F", X"AF", X"47", X"6F", --3DD0
  X"67", X"3A", X"6E", X"73", X"5F", X"3E", X"BF", X"93", --3DD8
  X"E6", X"F8", X"6F", X"CB", X"15", X"CB", X"14", X"AF", --3DE0
  X"CB", X"15", X"CB", X"14", X"09", X"22", X"86", X"7B", --3DE8
  X"01", X"00", X"58", X"09", X"3E", X"62", X"77", X"23", --3DF0
  X"77", X"23", X"77", X"C9", X"2B", X"3A", X"79", X"7B", --3DF8
  X"CB", X"4F", X"28", X"03", X"23", X"23", X"23", X"3A", --3E00
  X"82", X"7B", X"4F", X"0D", X"0D", X"3E", X"62", X"77", --3E08
  X"23", X"3A", X"79", X"7B", X"CB", X"4F", X"20", X"02", --3E10
  X"2B", X"2B", X"0D", X"20", X"F0", X"C9", X"3A", X"79", --3E18
  X"7B", X"CB", X"4F", X"20", X"11", X"3A", X"6F", X"73", --3E20
  X"CB", X"57", X"20", X"05", X"21", X"69", X"7E", X"18", --3E28
  X"14", X"21", X"79", X"7E", X"18", X"0F", X"3A", X"6F", --3E30
  X"73", X"CB", X"57", X"20", X"05", X"21", X"49", X"7E", --3E38
  X"18", X"03", X"21", X"59", X"7E", X"22", X"80", X"7B", --3E40
  X"C9", X"00", X"05", X"1F", X"FA", X"2F", X"FF", X"4F", --3E48
  X"FA", X"4C", X"78", X"92", X"14", X"11", X"22", X"10", --3E50
  X"A1", X"00", X"05", X"1F", X"FA", X"2F", X"FF", X"2F", --3E58
  X"FA", X"4C", X"78", X"4A", X"12", X"09", X"12", X"05", --3E60
  X"0A", X"A0", X"00", X"5F", X"F8", X"FF", X"F4", X"5F", --3E68
  X"F2", X"1E", X"32", X"28", X"49", X"44", X"88", X"85", --3E70
  X"08", X"A0", X"00", X"5F", X"F8", X"FF", X"F4", X"5F", --3E78
  X"F2", X"1E", X"32", X"28", X"51", X"48", X"90", X"50", --3E80
  X"A0", X"01", X"78", X"02", X"58", X"02", X"00", X"00", --3E88
  X"00", X"10", X"B0", X"02", X"90", X"03", X"00", X"00", --3E90
  X"00", X"60", X"88", X"00", X"70", X"01", X"00", X"00", --3E98
  X"00", X"60", X"50", X"02", X"50", X"04", X"00", X"00", --3EA0
  X"00", X"A0", X"88", X"00", X"50", X"02", X"00", X"00", --3EA8
  X"00", X"A0", X"88", X"02", X"60", X"04", X"00", X"00", --3EB0
  X"00", X"F0", X"90", X"00", X"58", X"03", X"00", X"00", --3EB8
  X"00", X"98", X"48", X"00", X"40", X"02", X"00", X"00", --3EC0
  X"00", X"01", X"78", X"02", X"38", X"02", X"00", X"00", --3EC8
  X"00", X"38", X"B0", X"02", X"40", X"04", X"00", X"00", --3ED0
  X"00", X"28", X"90", X"00", X"38", X"01", X"00", X"00", --3ED8
  X"00", X"28", X"78", X"02", X"30", X"03", X"00", X"00", --3EE0
  X"00", X"48", X"80", X"00", X"30", X"02", X"00", X"00", --3EE8
  X"00", X"70", X"70", X"02", X"30", X"05", X"00", X"00", --3EF0
  X"00", X"68", X"B0", X"00", X"40", X"01", X"00", X"00", --3EF8
  X"00", X"68", X"98", X"02", X"38", X"05", X"00", X"00", --3F00
  X"00", X"90", X"98", X"02", X"38", X"06", X"00", X"00", --3F08
  X"00", X"90", X"70", X"00", X"30", X"03", X"00", X"00", --3F10
  X"00", X"B8", X"A0", X"00", X"60", X"04", X"00", X"00", --3F18
  X"00", X"C0", X"98", X"02", X"40", X"08", X"00", X"00", --3F20
  X"00", X"B8", X"50", X"00", X"38", X"05", X"00", X"00", --3F28
  X"00", X"C8", X"78", X"02", X"38", X"08", X"00", X"00", --3F30
  X"00", X"F0", X"98", X"00", X"40", X"06", X"00", X"00", --3F38
  X"00", X"F0", X"70", X"00", X"38", X"07", X"00", X"00", --3F40
  X"00", X"ED", X"4B", X"86", X"7B", X"21", X"00", X"58", --3F48
  X"09", X"EB", X"21", X"30", X"75", X"09", X"01", X"03", --3F50
  X"00", X"ED", X"B0", X"C9", X"00", X"ED", X"B0", X"C9", --3F58
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3F60
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3F68
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3F70
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3F78
  X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"80", --3F80
  X"00", X"11", X"00", X"58", X"21", X"24", X"5F", X"ED", --3F88
  X"B0", X"C9", X"01", X"80", X"00", X"11", X"85", X"58", --3F90
  X"21", X"24", X"5F", X"7E", X"3C", X"3D", X"20", X"02", --3F98
  X"3E", X"64", X"CB", X"F7", X"12", X"23", X"13", X"0D", --3FA0
  X"20", X"F1", X"C9", X"21", X"80", X"58", X"0E", X"80", --3FA8
  X"3E", X"42", X"77", X"23", X"0D", X"20", X"FB", X"0E", --3FB0
  X"FF", X"77", X"23", X"0D", X"00", X"00", X"00", X"00", --3FB8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3FC0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3FC8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3FD0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3FD8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3FE0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3FE8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3FF0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00");--3FF8

begin

  process (clk)
  begin
    if(rising_edge(clk)) then
      if wr='1' then
        ram(to_integer(unsigned(addr))) <= din;
      end if;
      dout <= ram(to_integer(unsigned(addr)));
    end if; 
  end process;

end behavioral;
