library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library UNISIM;
use UNISIM.vcomponents.all;

entity vram is port(
    clk     : in  std_logic
  ; rd      : in  std_logic
  ; wr      : in  std_logic
  ; addr    : in  std_logic_vector(13 downto 0)
  ; dataout : out std_logic_vector( 7 downto 0)
);
end vram;

architecture Behavioral of vram is

type EN_a is array(7 downto 0) of std_logic;
type Arr_d is array(7 downto 0) of std_logic_vector(7 downto 0);
signal ENA : EN_a;
signal DOA : Arr_d;

begin

    process(addr, rd, DOA)
    variable i : integer;
    begin
        dataout <= (others => '0');
        for i in 0 to 7 loop
            ENA(i) <= '0';
            if (rd='1' and to_integer(unsigned(addr(13 downto 11))) = i) then
                ENA(i) <= '1';
                dataout <= DOA(i);
            end if;
        end loop;
    end process;

  ram0 : RAMB16_S9
  generic map (
      write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    , INIT_00   => X"9898989898989898989898989898989898989898989898989898989898989898"
    , INIT_01   => X"9898000000000000000000ffffffffffff0000ff0000ff000000000000009898"
    , INIT_02   => X"9898e0ffff03ff8feaff07000000000000fc7f00c0ff01fc7fe001fc03009898"
    , INIT_03   => X"989800f4ffff0300000000000000000000000f00000000000000fcffff009898"
    , INIT_04   => X"989800f9ff000000000000000000000000000000000000000000e0ff0f039898"
    , INIT_05   => X"9898007f0000000000000000000000000000000000f8fffffffffff03f009898"
    , INIT_06   => X"98983000000080ff68471c0000000000000000000000000000fe0100fe019898"
    , INIT_07   => X"989800437e003c3c001f3f7c1e7e1e9f071f3f7efc1ff83fc03f0000c0079898"
    , INIT_08   => X"6262626262626262626262626262626262626262626262626262626262626262"
    , INIT_09   => X"6262000000000000000080ffffffffffff0000ff0000ff000000000000006262"
    , INIT_0a   => X"6262f0ffff83ff0305ff03000000000000f07f00807f00f87fc003fc07006262"
    , INIT_0b   => X"626200e8ffff0100000000000000000000000600000000000000f8ffff016262"
    , INIT_0c   => X"626200fe7f000000000000000000000000000000000000000000f8ff0f076262"
    , INIT_0d   => X"6262801f0000000000000000000000000000000000f8ffffffff7fe07f006262"
    , INIT_0e   => X"6262c0010000f87ffc7f0e6002300020007680370000000000fe0100fc016262"
    , INIT_0f   => X"6262c000f0003c38001f7f7c1e7f1c9e071e3e3ebc1ffc7fc03f000080076262"
    , INIT_10   => X"1616161616161616161616161616161616161616161616161616161616161616"
    , INIT_11   => X"1616000000000000000080ffffffffffff0000ff0000ff000000000000001616"
    , INIT_12   => X"1616f8ffffc7ff0100fc00000000000000e07f00001f00e03fc007fe0f001616"
    , INIT_13   => X"161600d0ffff0000000000000000000000000200000000000000f8ffff011616"
    , INIT_14   => X"161600fd3f00000000000000000000000000000000400f00c001feff0f041616"
    , INIT_15   => X"1616800f0000000000000000000000000000000000f0ffffffff1fe07f001616"
    , INIT_16   => X"1616000f0000f87ffe7f0e3803703e38e17fd03fd833000700ff0100fc011616"
    , INIT_17   => X"1616300080017c18003f3e3e9e3f1c9e071e1f3e1e3efcffc03f000080071616"
    , INIT_18   => X"bcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbc"
    , INIT_19   => X"bcbc000000000000000000ffffffff0fff0100ff0000ff00000c00000000bcbc"
    , INIT_1a   => X"bcbcfcffffe7ff00003000000000000000c07f00000400c03f800fff1f00bcbc"
    , INIT_1b   => X"bcbc00e8ff3f0000000000000000000000000000000000000000f0ffff01bcbc"
    , INIT_1c   => X"bcbc80fc1f00000000000000000000000000000000e0dff5f88bfffe1f00bcbc"
    , INIT_1d   => X"bcbc80070000000000000000000000000000000000f081ffefff07c07f00bcbc"
    , INIT_1e   => X"bcbc007f0000fc7ffc3f1c3c0ff83cbeff3ff87ff87f801f00ff0000f803bcbc"
    , INIT_1f   => X"bcbc080000007c1cc03fbc1f9c7f1e0e073f1f3e1e3cfcffc03f00000007bcbc"
    , INIT_20   => X"a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3"
    , INIT_21   => X"a3a3000000000000000000c3ffffff00fc00c0ff0100ff00001a00000000a3a3"
    , INIT_22   => X"a3a3e4ffffff7f00000000000000000000c07f00000000801f009fff3f00a3a3"
    , INIT_23   => X"a3a300f4ff1f0000000000000000000000000000000000000000e0ffef01a3a3"
    , INIT_24   => X"a3a300ff0700000000000000000000000000000000e0fffffffffffd1f00a3a3"
    , INIT_25   => X"a3a3c00300000000000000000000000000000000008001d600ff0180ff00a3a3"
    , INIT_26   => X"a3a300ff0100fe3ffe3f1e3c0ff83c0eff3ffc7ff83fc00f007f0000f003a3a3"
    , INIT_27   => X"a3a338000000f83cc03f8c1f1e7f3e1e073e1c1e1c7c7e7fc07f0000000aa3a3"
    , INIT_28   => X"0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d"
    , INIT_29   => X"0d0d00feff0100000000c002f0ff0700f00040c10600bf00003c000000000d0d"
    , INIT_2a   => X"0d0d28ffffff3f00000000000000000000803f00000000000f00bfff7f000d0d"
    , INIT_2b   => X"0d0d00f8ff0f0000000000000000000000000000000000000000e0ffcf030d0d"
    , INIT_2c   => X"0d0d80fe0300000000000000000000000000000000f8ffffffffffff1f000d0d"
    , INIT_2d   => X"0d0dc001000000000000000000000000000000000000000000fe0080ff000d0d"
    , INIT_2e   => X"0d0d00ff0700fc3efe3f1e1c1f7c3c0eff3ffe7ff83fe01f807f0000f0030d0d"
    , INIT_2f   => X"0d0d70000000f07de01fce3f9e7f3c1e1e3e1c1e0c7c3efcc0ff0000000a0d0d"
    , INIT_30   => X"6161616161616161616161616161616161616161616161616161616161616161"
    , INIT_31   => X"616100ffff01fc7f06002001007c0000c000404208000f01007a000000006161"
    , INIT_32   => X"616150fdffff0f00000000000000000000801f00000000000e00feffff006161"
    , INIT_33   => X"616100f4ff070000000000000000000000000000000000000000c0ff8f036161"
    , INIT_34   => X"616100ff0100000000000000000000000000000000f8fffffffffffd3f006161"
    , INIT_35   => X"616140000000000000000000000000000000000000000000007e0000ff006161"
    , INIT_36   => X"616100ff0f007e1cfa1f1e1c0e7e3e1cff3fff3ffe1ff03f807f0000e0036161"
    , INIT_37   => X"6161f0000000f07ff01fcf3fdfff3e1c3c7e3e1e0c1e1ef880ff0000000c6161"
    , INIT_38   => X"3232323232323232323232323232323232323232323232323232323232323232"
    , INIT_39   => X"323200ffff03fe1f1800180000000000000340003200030200f4007800003232"
    , INIT_3a   => X"323280faffff0700000000000000000000000f00000000000400feffff003232"
    , INIT_3b   => X"323200faff030000000000000000000000000000000000000000c0ff8f033232"
    , INIT_3c   => X"323200ff0000000000000000000000000000000000f0fffffffffffa3f003232"
    , INIT_3d   => X"32322000000080e10000000000000000000000000000000000fe0000ff013232"
    , INIT_3e   => X"323200cf1f003e1c801f1e3c1c3e1e0f3f1efe7ffc1ff83f803f0000e0073232"
    , INIT_3f   => X"3232e0030000803ff01fff3fdf3f0e1e7c7e3e1e1c1e1ff801ff0100000c3232"
  )
  port map (
      DI    => "00000000"
    , DIP   => "0"
    , DO    => DOA(0)
    , ADDR  => addr(10 downto 0)
    , CLK   => clk
    , EN    => ENA(0)
    , WE    => wr
    , SSR   => '0'
  );

  ram1 : RAMB16_S9
  generic map (
      write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    , INIT_00   => X"9898e0070000807ff01ffe1ffe3f0e0ef07f3e3f1e1e3ef001ff010000f89898"
    , INIT_01   => X"989800ff3f001f1edc3f0f7f3f38fe1ffe3efc071f7ef03f80ff000000f09898"
    , INIT_02   => X"989800e0ffff0100000000000000000000000000000000000000000000e09898"
    , INIT_03   => X"98980000fcffff0f0000000000000000000000000000000000c0800000ff9898"
    , INIT_04   => X"9898000080ffffff7f0000000000000000000000020000bcff3c020100f09898"
    , INIT_05   => X"9898000000f8ffffffff070000000000102104080f0000ffffff530000f89898"
    , INIT_06   => X"9898000000f8ffefffffff3f00000001000000000000ea00fe1f871a00509898"
    , INIT_07   => X"9898000000f03f00000000f0ff0100000000000000f0400041bff000a03e9898"
    , INIT_08   => X"6262e01f0000f07fc01fff3dfe731e0ef03f3c3f3f1f7ef800fe010000f06262"
    , INIT_09   => X"626200feff001f1efc1f0f7f3e38fc0f3f3ef8871f3ef81f807f000000f86262"
    , INIT_0a   => X"626200c0ffff0700000000000000000000000000000000000060000000f06262"
    , INIT_0b   => X"62620000f8ffff3f0000000000000000000000000000000000d8800000fe6262"
    , INIT_0c   => X"6262000080ffffffff01000000000000840003000200c0427f42040100f86262"
    , INIT_0d   => X"6262000000f8ffffffff0f00001ce38e13210410008000fff7fea30000f06262"
    , INIT_0e   => X"6262000000f8ffc7ffc0ff7f0000000100000000000050000000831400686262"
    , INIT_0f   => X"6262000000f07f00000000f0ff0300000000000000f0200000bff800503f6262"
    , INIT_10   => X"1616c03f0000f03f003eff3cfe733e0ef03f3e0fff1ffefc00fe010000f01616"
    , INIT_11   => X"161600feff011e1efc0f0f7f1e78fc0f7e3ef00f0f3ef00f007f000000f81616"
    , INIT_12   => X"161600c0ffff0f000000000000000000000000000000000000c0010000fc1616"
    , INIT_13   => X"16160000f8ffff7f0000000000000000000000000000000000f8000000f81616"
    , INIT_14   => X"1616000000ffffffff0300000000000088c002000400e08f1cf1050000f81616"
    , INIT_15   => X"1616000000f8ffffffff1f0000a0949024420420008000ffffffa70000f01616"
    , INIT_16   => X"1616000000f8ff077f80ffff000000010000000000008e010000802f00741616"
    , INIT_17   => X"1616000000f0ff00000000e0ff0f00000000000000f8200000bff800b03f1616"
    , INIT_18   => X"bcbcc07f0000f03f003e7e1cfe703e0cf83f3e3fff1fffff01fe010000e0bcbc"
    , INIT_19   => X"bcbc00fcff03078cff1f033e0ff8fc1f0f7ef08f0f3cf007007e000000fcbcbc"
    , INIT_1a   => X"bcbc0080ffff1f000000000000000000000000000000000000c0070000febcbc"
    , INIT_1b   => X"bcbc0000f0ffffff0100000000000000000000000000000000a8000000f0bcbc"
    , INIT_1c   => X"bcbc000000ffffffff0f00000000000088200200040050bd42bd0a0000f8bcbc"
    , INIT_1d   => X"bcbc000000f8ffffffff7f00002097902442044000c0007ff883470100e0bcbc"
    , INIT_1e   => X"bcbc000000f8ff037e80ffff030000020000000000003f0f00f0802f003abcbc"
    , INIT_1f   => X"bcbc000000e0ff01000000e0ff1f00000000000000f8500000bf7d00d81fbcbc"
    , INIT_20   => X"a3a380ff0100fe7f001e7e1c7f303e0ef83f3e9fff1ffeff00fe010000c0a3a3"
    , INIT_21   => X"a3a300fcff0f031c87bf033c0ff8fc1f0f74f08f0f38c003007e000000fca3a3"
    , INIT_22   => X"a3a30080ffff7f000000000000000000000000000000000000c00f0000ffa3a3"
    , INIT_23   => X"a3a30000e0ffffff0300000000000000000000000000000000ac000000e0a3a3"
    , INIT_24   => X"a3a3000000feffffff1f00000000000088200200040058fe24ff160000fca3a3"
    , INIT_25   => X"a3a3000000f8ffffffffff00002094902482048010c00c1fe000820700e0a3a3"
    , INIT_26   => X"a3a3000000f8ff013c00fffd07000000000000000080fff0ffcfc053003da3a3"
    , INIT_27   => X"a3a3000000e0ff03000000c0ff3f00000000000000fc280000bf7f00f41fa3a3"
    , INIT_28   => X"0d0d80ff0300fe3f001f7f3c3f703c0eff1f3e0fff1ffc7f00fe010000e00d0d"
    , INIT_29   => X"0d0d00f8ff1f001c009f0330022000100000000000780000003c000000f80d0d"
    , INIT_2a   => X"0d0d0000ffffff000000000000000000000000000000000000801f0080ff0d0d"
    , INIT_2b   => X"0d0d0000e0ffffff07000000000000000000000000000000005f000100e00d0d"
    , INIT_2c   => X"0d0d000000feffffff3f000000000000881002220b005c9c0039120000fc0d0d"
    , INIT_2d   => X"0d0d000000f8ffffffffff0100a1e35023120700138070070000c00e00c00d0d"
    , INIT_2e   => X"0d0d000000f8ff00100000fc1f0000000000000000c0ff000080c063003a0d0d"
    , INIT_2f   => X"0d0d000000e0ffc7010000c0ffff00000000000000fc180000bf3f00fa1f0d0d"
    , INIT_30   => X"616180ff07007e7e001f1f3e3f787c1fff3efc0f3f3ff83f00ff010000e06161"
    , INIT_31   => X"616100f0ff7f000000000000000000000000000000000000003c000000e06161"
    , INIT_32   => X"61610000feffff030000000000000000000000000000000000803f00c0ff6161"
    , INIT_33   => X"61610000c0ffffff1f0000000000000000000000000000000041180100f06161"
    , INIT_34   => X"6161000000fcffffffff000000000000101102920800e66100862b0000fc6161"
    , INIT_35   => X"6161000000f8ffffffffff0700008000000000000c8081000000800f00e06161"
    , INIT_36   => X"6161000000f0ff00000000f83f0000000000000000c0ff400081e001803d6161"
    , INIT_37   => X"616100000080ffbf000000c0ffff01000000000000fe240000df3f00f51f6161"
    , INIT_38   => X"323200ff1f003f1e001f0e7f3f78fe1f7e1efc0f1f7ef83f00ff000000f03232"
    , INIT_39   => X"323200f0ffff0000000000000000000000000000000000000018000000c03232"
    , INIT_3a   => X"32320000feffff070000000000000000000000000000000000803f0080ff3232"
    , INIT_3b   => X"32320000c0ffffff3f00000000000000000000000200003c007e7e0100f03232"
    , INIT_3c   => X"3232000000fcffffffff010000000000f01104940800ff3e007c510000f83232"
    , INIT_3d   => X"3232000000f8ffffffffff0f0000000100000000000002070000041f00e03232"
    , INIT_3e   => X"3232000000f07f00000000f87f0000000000000000e0ff808020e001403f3232"
    , INIT_3f   => X"323200000000fc7f000000c0ffff03000000000000ff1600009f1f00fb0f3232"
  )
  port map (
      DI    => "00000000"
    , DIP   => "0"
    , DO    => DOA(1)
    , ADDR  => addr(10 downto 0)
    , CLK   => clk
    , EN    => ENA(1)
    , WE    => wr
    , SSR   => '0'
  );

  ram2 : RAMB16_S9
  generic map (
      write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    , INIT_00   => X"989800000000f03f000000c0ffff0f000000000080000b00420f0f80fd079898"
    , INIT_01   => X"9898000000000000000000000000fcff00000000ffaf0000e00000f57f009898"
    , INIT_02   => X"9898000000000000000000000000e0ffff030070000100000000f4ffff019898"
    , INIT_03   => X"989800fc3f0000000000000000000000f8ff1f085f550207375007c07f009898"
    , INIT_04   => X"9898ffffffffdcf7ffff77dffd7f00e0ffffe0ffff03c003a0fe7f0018009898"
    , INIT_05   => X"9898fc3ffc3f505495e477dbc17e000000000000e0af45adfe001f0000009898"
    , INIT_06   => X"9898989898989898989898989898989898989898989898989898989898989898"
    , INIT_07   => X"9898989898989898989898989898989898989898989898989898989898989898"
    , INIT_08   => X"626200000000801f000000c0ffff1f0000000000c08007f881000640ff016262"
    , INIT_09   => X"6262000000000000000000000000f8ff010000007f1f003ff00000fb7f006262"
    , INIT_0a   => X"6262000000000000000000000000c0ffff070078000100000c00faffff016262"
    , INIT_0b   => X"626200e00f00700f0000700000000000f8ff3f04afa001030ae807807e006262"
    , INIT_0c   => X"6262fc3ffc3f501400007000000000f8ffffc0ffff00e00160ff7f0018006262"
    , INIT_0d   => X"6262e007e007505455e276dbc16e000000000000c05f877d3f001e0000006262"
    , INIT_0e   => X"6262626262626262626262626262626262626262626262626262626262626262"
    , INIT_0f   => X"6262626262626262626262626262626262626262626262626262626262626262"
    , INIT_10   => X"161600000000000c000000c09fff7f0000000000c0c00b00000700a0ff001616"
    , INIT_11   => X"1616ce24894ccecea8a9b0ab9324fcff030000803f07e0c0ff0080fd7f001616"
    , INIT_12   => X"161600000000004024764462236680ffff1f007c000100200300f4ffff011616"
    , INIT_13   => X"16160080010050110000700000000000f8ffff005750008103f40f007f001616"
    , INIT_14   => X"1616e007e007501400007000000000feff7f80ff3e00f800b0ff3f0010001616"
    , INIT_15   => X"161680018001505455e176dbc16e00000000000000bf04aa0f00180000001616"
    , INIT_16   => X"1616161616161616161616161616161616161616161616161616161616161616"
    , INIT_17   => X"1616161616161616161616161616161616161616161616161616161616161616"
    , INIT_18   => X"bcbc000000000000000000c001ffff0000000000e0f00500000300507f00bcbc"
    , INIT_19   => X"bcbc28a5daaaa8a828aa282aa954f8ff070000c01f031800f00040ff7f00bcbc"
    , INIT_1a   => X"bcbc0000000000c056456c55545500fffb3e0036000200d40080fbffff01bcbc"
    , INIT_1b   => X"bcbc0000000050170000700000000000f8ffff010ba8004100ea1f007f00bcbc"
    , INIT_1c   => X"bcbc800180015014c7c773ceb93c00ffff3f00801d007c00e8ff3f000000bcbc"
    , INIT_1d   => X"bcbc000000005c5452ef76dfc16e000000000000005c03f4030010000000bcbc"
    , INIT_1e   => X"bcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbc"
    , INIT_1f   => X"acbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbcbc"
    , INIT_20   => X"a3a30000000000000000000000fcff0100000000f0f80200110100b01f00a3a3"
    , INIT_21   => X"a3a308b5aaaaa8a828aa282aa956fcff0f0000c00f0304000000a0ffff00a3a3"
    , INIT_22   => X"a3a300800100004055455455545500fef8ff002b8003802a00c0f5feff00a3a3"
    , INIT_23   => X"a3a30000000050140000700000000000f8ffff0707d000a000f61f003e00a3a3"
    , INIT_24   => X"a3a300000000509448e877dffd7e0000000000002e002b00f4ff3f000000a3a3"
    , INIT_25   => X"a3a300000000449448e877dfc17e00000000000000e80338000000000000a3a3"
    , INIT_26   => X"a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3"
    , INIT_27   => X"ffa3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3"
    , INIT_28   => X"0d0d0000000000000000000000f8ff0700000000f87c0180100000d81f000d0d"
    , INIT_29   => X"0d0d0cad8bacccccb8ea303ba975f8ff3f0000e007010000001f50ffff000d0d"
    , INIT_2a   => X"0d0d00e007000040546644675566007ef8ff81354006501500753afcff000d0d"
    , INIT_2b   => X"0d0d80018001dcf7ffff77dffd7f0000f8ffff0f01e800c000fb3f003e000d0d"
    , INIT_2c   => X"0d0d000000005054d26b76dfcd6600000000000015803500eaff3f0000000d0d"
    , INIT_2d   => X"0d0d000000007c1c876f73cec136000000000000008003080000000000000d0d"
    , INIT_2e   => X"0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d"
    , INIT_2f   => X"e00e0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d0d"
    , INIT_30   => X"61610000000000000000000000f0ff0f00000000fcbe0240a00000f43f006161"
    , INIT_31   => X"616128a58aaaa888a8aa282aa954f0ff7f0000e001010000007fb0ffff006161"
    , INIT_32   => X"616100fc3f00cc4c544544555545003cf8ff8336801da80f80bc0df8ff006161"
    , INIT_33   => X"6161e007e0070400000074d105400000fefffb1f00f080e080fe3f003c006161"
    , INIT_34   => X"616100000000505415ea70dbc10e0000000000002ac01a00f6ef3f0000006161"
    , INIT_35   => X"6161000000000000000000000000000000000000000000000000000000006161"
    , INIT_36   => X"6161616161616161616161616161616161616161616161616161616161616161"
    , INIT_37   => X"ea62616161616161616161616161616161616161616161616161616161616161"
    , INIT_38   => X"3232000000000000000000000000ff3f00000000fe5e0100c00000fa3f003232"
    , INIT_39   => X"3232cea48a4aa88ea8a9a82b9154e0ffff0100f00001000000ffd8ffff003232"
    , INIT_3a   => X"323200ffff00cc4c2445445523450008f8ff0f1b60eaff07505f02e0ff003232"
    , INIT_3b   => X"3232fc3ffc3f0400000074d105400080fffff17f00f880f840fd7f003c003232"
    , INIT_3c   => X"323200000000505415e973dbc13e00000000000055012b087b833f0000003232"
    , INIT_3d   => X"3232000000000000000000000000000000000000000000000000000000003232"
    , INIT_3e   => X"3232323232323232323232323232323232323232323232323232323232323232"
    , INIT_3f   => X"2a32323232323232323232323232323232323232323232323232323232323232"
  )
  port map (
      DI    => "00000000"
    , DIP   => "0"
    , DO    => DOA(2)
    , ADDR  => addr(10 downto 0)
    , CLK   => clk
    , EN    => ENA(2)
    , WE    => wr
    , SSR   => '0'
  );

  ram3 : RAMB16_S9
  generic map (
      write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    , INIT_00   => X"7878787878787878787878787878787878787878787878787878787878787878"
    , INIT_01   => X"78780a0a0a0a0a0a090a09010101010101090901090a01090a0a0a0a0a0a7878"
    , INIT_02   => X"78380a0a0a0a02010101010202020202020101020101010101020a0a0a0a7878"
    , INIT_03   => X"78380a0a0a020202020202020202020202020102020202020202020a0a0a7878"
    , INIT_04   => X"78380a0a0202020202020202020202020202020202464646464646320a0a7878"
    , INIT_05   => X"78380a020202060602020202020202020202020202464646464646020a0a7878"
    , INIT_06   => X"78380901010246464646464646464646464646464646464606460602020a7878"
    , INIT_07   => X"78380901010146464646464646464646464646464646464646460602020a7878"
    , INIT_08   => X"78380a0202064646464646464646464646464646464646460646460202017878"
    , INIT_09   => X"78380a0a0a024646464646464646464646464646464646464646020202017878"
    , INIT_0a   => X"78380a0a0a0a0202020202020202424242424242420202020343434301017878"
    , INIT_0b   => X"78380a0a0a0a0a02020202020202424242424242420203040343580302017878"
    , INIT_0c   => X"78380a0a0a0a0a0a0a0202020202424245454542420304202084044302017878"
    , INIT_0d   => X"78380a0a0a0a0a0a0a0a020202454545454545424204200c0c0c040402017878"
    , INIT_0e   => X"78380a0a0a0a0a0a0a0a0a0a02024245424242424204042020200404020a7878"
    , INIT_0f   => X"78380a0a0a0a0a0a0a0a0a0a0a020202020202020204202020040403020a7878"
    , INIT_10   => X"78380a0a0a0a0a0a0a0a0a0a0a0a02020202020204202020200444020a0a7878"
    , INIT_11   => X"78384747474747474747474747470a0a0202020404202020200402020a0a7878"
    , INIT_12   => X"78384641414647474747474747470a0a0a0202040420202020200a0a0a0a7878"
    , INIT_13   => X"78384121514147474747474747470a0a0a0a02022020042004020a0a0a0a7878"
    , INIT_14   => X"78382151215147474747474747470a0a0a0a0a0a04040404020a0a0a0a0a7878"
    , INIT_15   => X"78380442044247474747474747470a0a0a0a0a0a0a0a0a0a0a0a0a0a0a0a7878"
    , INIT_16   => X"7838383838383838383838383838383838383838383838383838383838787878"
    , INIT_17   => X"7878787878787878787878787878787878787878787878787878787878787878"
  )
  port map (
      DI    => "00000000"
    , DIP   => "0"
    , DO    => DOA(3)
    , ADDR  => addr(10 downto 0)
    , CLK   => clk
    , EN    => ENA(3)
    , WE    => wr
    , SSR   => '0'
  );

    RAMB : for i in 4 to 7 generate
    RAMB16_S9_inst : RAMB16_S9
    generic map (
        write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    )
    port map (
        DO => DOA(i),      -- 8-bit Data Output
        ADDR => addr(10 downto 0),  -- 11-bit Address Input
        CLK => clk,    -- Clock
        DI => "00000000",      -- 8-bit Data Input
        DIP => "0",
        EN => ENA(i),      -- RAM Enable Input
        SSR => '0',    -- Synchronous Set/Reset Input
        WE => wr       -- Write Enable Input
    );
    end generate;

--  ram4 : RAMB16_S9
--  generic map (
--      write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
--  )
--  port map (
--      DI    => "00000000"
--    , DO    => dataout
--    , ADDR  => "00000000000"
--    , CLK   => clk
--    , EN    => ram4en
--    , WE    => '0'
--    , SSR   => '0'
--  );

end Behavioral;
