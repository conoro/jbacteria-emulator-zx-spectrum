library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is port(
    clk   : in  std_logic;
    addr  : in  std_logic_vector(9 downto 0);
    dout  : out std_logic_vector(7 downto 0));
end rom;

architecture behavioral of rom is

  type rom_t is array (0 to 1023) of std_logic_vector(7 downto 0);
  signal rom : rom_t := (
  X"F3", X"31", X"40", X"7C", X"C3", X"F6", X"64", X"11", --0000
  X"2A", X"5D", X"5C", X"22", X"5F", X"5C", X"18", X"43", --0008
  X"C3", X"F2", X"15", X"FF", X"FF", X"FF", X"FF", X"FF", --0010
  X"2A", X"5D", X"5C", X"7E", X"CD", X"7D", X"00", X"D0", --0018
  X"CD", X"74", X"00", X"18", X"F7", X"FF", X"FF", X"FF", --0020
  X"C3", X"5B", X"33", X"FF", X"FF", X"FF", X"FF", X"FF", --0028
  X"C5", X"2A", X"61", X"5C", X"E5", X"C3", X"9E", X"16", --0030
  X"F5", X"E5", X"2A", X"78", X"5C", X"23", X"22", X"78", --0038
  X"5C", X"7C", X"B5", X"20", X"03", X"FD", X"34", X"40", --0040
  X"C5", X"D5", X"CD", X"BF", X"02", X"D1", X"C1", X"E1", --0048
  X"F1", X"FB", X"C9", X"E1", X"6E", X"FD", X"75", X"00", --0050
  X"ED", X"7B", X"3D", X"5C", X"C3", X"C5", X"16", X"FF", --0058
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F5", X"E5", --0060
  X"2A", X"B0", X"5C", X"7C", X"B5", X"20", X"01", X"E9", --0068
  X"E1", X"F1", X"ED", X"45", X"2A", X"5D", X"5C", X"23", --0070
  X"22", X"5D", X"5C", X"7E", X"C9", X"FE", X"21", X"D0", --0078
  X"FE", X"0D", X"C8", X"FE", X"10", X"D8", X"FE", X"18", --0080
  X"3F", X"D8", X"23", X"FE", X"16", X"38", X"01", X"23", --0088
  X"37", X"22", X"5D", X"5C", X"C9", X"BF", X"52", X"4E", --0090
  X"C4", X"49", X"4E", X"4B", X"45", X"59", X"A4", X"50", --0098
  X"C9", X"46", X"CE", X"50", X"4F", X"49", X"4E", X"D4", --00A0
  X"53", X"43", X"52", X"45", X"45", X"4E", X"A4", X"41", --00A8
  X"54", X"54", X"D2", X"41", X"D4", X"54", X"41", X"C2", --00B0
  X"56", X"41", X"4C", X"A4", X"43", X"4F", X"44", X"C5", --00B8
  X"56", X"41", X"CC", X"4C", X"45", X"CE", X"53", X"49", --00C0
  X"CE", X"43", X"4F", X"D3", X"54", X"41", X"CE", X"41", --00C8
  X"53", X"CE", X"41", X"43", X"D3", X"41", X"54", X"CE", --00D0
  X"4C", X"CE", X"45", X"58", X"D0", X"49", X"4E", X"D4", --00D8
  X"53", X"51", X"D2", X"53", X"47", X"CE", X"41", X"42", --00E0
  X"D3", X"50", X"45", X"45", X"CB", X"49", X"CE", X"55", --00E8
  X"53", X"D2", X"53", X"54", X"52", X"A4", X"43", X"48", --00F0
  X"52", X"A4", X"4E", X"4F", X"D4", X"42", X"49", X"CE", --00F8
  X"4F", X"D2", X"41", X"4E", X"C4", X"3C", X"BD", X"3E", --0100
  X"BD", X"3C", X"BE", X"4C", X"49", X"4E", X"C5", X"54", --0108
  X"48", X"45", X"CE", X"54", X"CF", X"53", X"54", X"45", --0110
  X"D0", X"44", X"45", X"46", X"20", X"46", X"CE", X"43", --0118
  X"41", X"D4", X"46", X"4F", X"52", X"4D", X"41", X"D4", --0120
  X"4D", X"4F", X"56", X"C5", X"45", X"52", X"41", X"53", --0128
  X"C5", X"4F", X"50", X"45", X"4E", X"20", X"A3", X"43", --0130
  X"4C", X"4F", X"53", X"45", X"20", X"A3", X"4D", X"45", --0138
  X"52", X"47", X"C5", X"56", X"45", X"52", X"49", X"46", --0140
  X"D9", X"42", X"45", X"45", X"D0", X"43", X"49", X"52", --0148
  X"43", X"4C", X"C5", X"49", X"4E", X"CB", X"50", X"41", --0150
  X"50", X"45", X"D2", X"46", X"4C", X"41", X"53", X"C8", --0158
  X"42", X"52", X"49", X"47", X"48", X"D4", X"49", X"4E", --0160
  X"56", X"45", X"52", X"53", X"C5", X"4F", X"56", X"45", --0168
  X"D2", X"4F", X"55", X"D4", X"4C", X"50", X"52", X"49", --0170
  X"4E", X"D4", X"4C", X"4C", X"49", X"53", X"D4", X"53", --0178
  X"54", X"4F", X"D0", X"52", X"45", X"41", X"C4", X"44", --0180
  X"41", X"54", X"C1", X"52", X"45", X"53", X"54", X"4F", --0188
  X"52", X"C5", X"4E", X"45", X"D7", X"42", X"4F", X"52", --0190
  X"44", X"45", X"D2", X"43", X"4F", X"4E", X"54", X"49", --0198
  X"4E", X"55", X"C5", X"44", X"49", X"CD", X"52", X"45", --01A0
  X"CD", X"46", X"4F", X"D2", X"47", X"4F", X"20", X"54", --01A8
  X"CF", X"47", X"4F", X"20", X"53", X"55", X"C2", X"49", --01B0
  X"4E", X"50", X"55", X"D4", X"4C", X"4F", X"41", X"C4", --01B8
  X"4C", X"49", X"53", X"D4", X"4C", X"45", X"D4", X"50", --01C0
  X"41", X"55", X"53", X"C5", X"4E", X"45", X"58", X"D4", --01C8
  X"50", X"4F", X"4B", X"C5", X"50", X"52", X"49", X"4E", --01D0
  X"D4", X"50", X"4C", X"4F", X"D4", X"52", X"55", X"CE", --01D8
  X"53", X"41", X"56", X"C5", X"52", X"41", X"4E", X"44", --01E0
  X"4F", X"4D", X"49", X"5A", X"C5", X"49", X"C6", X"43", --01E8
  X"4C", X"D3", X"44", X"52", X"41", X"D7", X"43", X"4C", --01F0
  X"45", X"41", X"D2", X"52", X"45", X"54", X"55", X"52", --01F8
  X"CE", X"43", X"4F", X"50", X"D9", X"42", X"48", X"59", --0200
  X"36", X"35", X"54", X"47", X"56", X"4E", X"4A", X"55", --0208
  X"37", X"34", X"52", X"46", X"43", X"4D", X"4B", X"49", --0210
  X"38", X"33", X"45", X"44", X"58", X"0E", X"4C", X"4F", --0218
  X"39", X"32", X"57", X"53", X"5A", X"20", X"0D", X"50", --0220
  X"30", X"31", X"51", X"41", X"E3", X"C4", X"E0", X"E4", --0228
  X"B4", X"BC", X"BD", X"BB", X"AF", X"B0", X"B1", X"C0", --0230
  X"A7", X"A6", X"BE", X"AD", X"B2", X"BA", X"E5", X"A5", --0238
  X"C2", X"E1", X"B3", X"B9", X"C1", X"B8", X"7E", X"DC", --0240
  X"DA", X"5C", X"B7", X"7B", X"7D", X"D8", X"BF", X"AE", --0248
  X"AA", X"AB", X"DD", X"DE", X"DF", X"7F", X"B5", X"D6", --0250
  X"7C", X"D5", X"5D", X"DB", X"B6", X"D9", X"5B", X"D7", --0258
  X"0C", X"07", X"06", X"04", X"05", X"08", X"0A", X"0B", --0260
  X"09", X"0F", X"E2", X"2A", X"3F", X"CD", X"C8", X"CC", --0268
  X"CB", X"5E", X"AC", X"2D", X"2B", X"3D", X"2E", X"2C", --0270
  X"3B", X"22", X"C7", X"3C", X"C3", X"3E", X"C5", X"2F", --0278
  X"C9", X"60", X"C6", X"3A", X"D0", X"CE", X"A8", X"CA", --0280
  X"D3", X"D4", X"D1", X"D2", X"A9", X"CF", X"2E", X"2F", --0288
  X"11", X"FF", X"FF", X"01", X"FE", X"FE", X"ED", X"78", --0290
  X"2F", X"E6", X"1F", X"28", X"0E", X"67", X"7D", X"14", --0298
  X"C0", X"D6", X"08", X"CB", X"3C", X"30", X"FA", X"53", --02A0
  X"5F", X"20", X"F4", X"2D", X"CB", X"00", X"38", X"E6", --02A8
  X"7A", X"3C", X"C8", X"FE", X"28", X"C8", X"FE", X"19", --02B0
  X"C8", X"7B", X"5A", X"57", X"FE", X"18", X"C9", X"CD", --02B8
  X"8E", X"02", X"C0", X"21", X"00", X"5C", X"CB", X"7E", --02C0
  X"20", X"07", X"23", X"35", X"2B", X"20", X"02", X"36", --02C8
  X"FF", X"7D", X"21", X"04", X"5C", X"BD", X"20", X"EE", --02D0
  X"CD", X"1E", X"03", X"D0", X"21", X"00", X"5C", X"BE", --02D8
  X"28", X"2E", X"EB", X"21", X"04", X"5C", X"BE", X"28", --02E0
  X"27", X"CB", X"7E", X"20", X"04", X"EB", X"CB", X"7E", --02E8
  X"C8", X"5F", X"77", X"23", X"36", X"05", X"23", X"3A", --02F0
  X"09", X"5C", X"77", X"23", X"FD", X"4E", X"07", X"FD", --02F8
  X"56", X"01", X"E5", X"CD", X"33", X"03", X"E1", X"77", --0300
  X"32", X"08", X"5C", X"FD", X"CB", X"01", X"EE", X"C9", --0308
  X"23", X"36", X"05", X"23", X"35", X"C0", X"3A", X"0A", --0310
  X"5C", X"77", X"23", X"7E", X"18", X"EA", X"42", X"16", --0318
  X"00", X"7B", X"FE", X"27", X"D0", X"FE", X"18", X"20", --0320
  X"03", X"CB", X"78", X"C0", X"21", X"05", X"02", X"19", --0328
  X"7E", X"37", X"C9", X"7B", X"FE", X"3A", X"38", X"2F", --0330
  X"0D", X"FA", X"4F", X"03", X"28", X"03", X"C6", X"4F", --0338
  X"C9", X"21", X"EB", X"01", X"04", X"28", X"03", X"21", --0340
  X"05", X"02", X"16", X"00", X"19", X"7E", X"C9", X"21", --0348
  X"29", X"02", X"CB", X"40", X"28", X"F4", X"CB", X"5A", --0350
  X"28", X"0A", X"FD", X"CB", X"30", X"5E", X"C0", X"04", --0358
  X"C0", X"C6", X"20", X"C9", X"C6", X"A5", X"C9", X"FE", --0360
  X"30", X"D8", X"0D", X"FA", X"9D", X"03", X"20", X"19", --0368
  X"21", X"54", X"02", X"CB", X"68", X"28", X"D3", X"FE", --0370
  X"38", X"30", X"07", X"D6", X"20", X"04", X"C8", X"C6", --0378
  X"08", X"C9", X"D6", X"36", X"04", X"C8", X"C6", X"FE", --0380
  X"C9", X"21", X"30", X"02", X"FE", X"39", X"28", X"BA", --0388
  X"FE", X"30", X"28", X"B6", X"E6", X"07", X"C6", X"80", --0390
  X"04", X"C8", X"EE", X"0F", X"C9", X"04", X"C8", X"CB", --0398
  X"68", X"21", X"30", X"02", X"20", X"A4", X"D6", X"10", --03A0
  X"FE", X"22", X"28", X"06", X"FE", X"20", X"C0", X"3E", --03A8
  X"5F", X"C9", X"3E", X"40", X"C9", X"F3", X"7D", X"CB", --03B0
  X"3D", X"CB", X"3D", X"2F", X"E6", X"03", X"4F", X"06", --03B8
  X"00", X"DD", X"21", X"D1", X"03", X"DD", X"09", X"3A", --03C0
  X"48", X"5C", X"E6", X"38", X"0F", X"0F", X"0F", X"F6", --03C8
  X"08", X"00", X"00", X"00", X"04", X"0C", X"0D", X"20", --03D0
  X"FD", X"0E", X"3F", X"05", X"C2", X"D6", X"03", X"EE", --03D8
  X"10", X"D3", X"FE", X"44", X"4F", X"CB", X"67", X"20", --03E0
  X"09", X"7A", X"B3", X"28", X"09", X"79", X"4D", X"1B", --03E8
  X"DD", X"E9", X"4D", X"0C", X"DD", X"E9", X"FB", X"C9", --03F0
  X"EF", X"31", X"27", X"C0", X"03", X"34", X"EC", X"6C");--03F8

begin

  process (clk)
  begin
    if rising_edge(clk) then
      dout <= rom(to_integer(unsigned(addr)));
    end if;
  end process;

end behavioral;
