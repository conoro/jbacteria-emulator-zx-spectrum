library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is port(
    clk   : in  std_logic;
    addr  : in  std_logic_vector(13 downto 0);
    dout  : out std_logic_vector(7 downto 0));
end rom;

architecture behavioral of rom is

  type rom_t is array (0 to 16383) of std_logic_vector(7 downto 0);
  signal rom : rom_t := (
  X"F3", X"AF", X"11", X"FF", X"FF", X"C3", X"CB", X"11", --0000
  X"2A", X"5D", X"5C", X"22", X"5F", X"5C", X"18", X"43", --0008
  X"C3", X"F2", X"15", X"FF", X"FF", X"FF", X"FF", X"FF", --0010
  X"2A", X"5D", X"5C", X"7E", X"CD", X"7D", X"00", X"D0", --0018
  X"CD", X"74", X"00", X"18", X"F7", X"FF", X"FF", X"FF", --0020
  X"C3", X"5B", X"33", X"FF", X"FF", X"FF", X"FF", X"FF", --0028
  X"C5", X"2A", X"61", X"5C", X"E5", X"C3", X"9E", X"16", --0030
  X"F5", X"E5", X"2A", X"78", X"5C", X"23", X"22", X"78", --0038
  X"5C", X"7C", X"B5", X"20", X"03", X"FD", X"34", X"40", --0040
  X"C5", X"D5", X"CD", X"BF", X"02", X"D1", X"C1", X"E1", --0048
  X"F1", X"FB", X"C9", X"E1", X"6E", X"FD", X"75", X"00", --0050
  X"ED", X"7B", X"3D", X"5C", X"C3", X"C5", X"16", X"FF", --0058
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F5", X"E5", --0060
  X"2A", X"B0", X"5C", X"7C", X"B5", X"20", X"01", X"E9", --0068
  X"E1", X"F1", X"ED", X"45", X"2A", X"5D", X"5C", X"23", --0070
  X"22", X"5D", X"5C", X"7E", X"C9", X"FE", X"21", X"D0", --0078
  X"FE", X"0D", X"C8", X"FE", X"10", X"D8", X"FE", X"18", --0080
  X"3F", X"D8", X"23", X"FE", X"16", X"38", X"01", X"23", --0088
  X"37", X"22", X"5D", X"5C", X"C9", X"BF", X"52", X"4E", --0090
  X"C4", X"49", X"4E", X"4B", X"45", X"59", X"A4", X"50", --0098
  X"C9", X"46", X"CE", X"50", X"4F", X"49", X"4E", X"D4", --00A0
  X"53", X"43", X"52", X"45", X"45", X"4E", X"A4", X"41", --00A8
  X"54", X"54", X"D2", X"41", X"D4", X"54", X"41", X"C2", --00B0
  X"56", X"41", X"4C", X"A4", X"43", X"4F", X"44", X"C5", --00B8
  X"56", X"41", X"CC", X"4C", X"45", X"CE", X"53", X"49", --00C0
  X"CE", X"43", X"4F", X"D3", X"54", X"41", X"CE", X"41", --00C8
  X"53", X"CE", X"41", X"43", X"D3", X"41", X"54", X"CE", --00D0
  X"4C", X"CE", X"45", X"58", X"D0", X"49", X"4E", X"D4", --00D8
  X"53", X"51", X"D2", X"53", X"47", X"CE", X"41", X"42", --00E0
  X"D3", X"50", X"45", X"45", X"CB", X"49", X"CE", X"55", --00E8
  X"53", X"D2", X"53", X"54", X"52", X"A4", X"43", X"48", --00F0
  X"52", X"A4", X"4E", X"4F", X"D4", X"42", X"49", X"CE", --00F8
  X"4F", X"D2", X"41", X"4E", X"C4", X"3C", X"BD", X"3E", --0100
  X"BD", X"3C", X"BE", X"4C", X"49", X"4E", X"C5", X"54", --0108
  X"48", X"45", X"CE", X"54", X"CF", X"53", X"54", X"45", --0110
  X"D0", X"44", X"45", X"46", X"20", X"46", X"CE", X"43", --0118
  X"41", X"D4", X"46", X"4F", X"52", X"4D", X"41", X"D4", --0120
  X"4D", X"4F", X"56", X"C5", X"45", X"52", X"41", X"53", --0128
  X"C5", X"4F", X"50", X"45", X"4E", X"20", X"A3", X"43", --0130
  X"4C", X"4F", X"53", X"45", X"20", X"A3", X"4D", X"45", --0138
  X"52", X"47", X"C5", X"56", X"45", X"52", X"49", X"46", --0140
  X"D9", X"42", X"45", X"45", X"D0", X"43", X"49", X"52", --0148
  X"43", X"4C", X"C5", X"49", X"4E", X"CB", X"50", X"41", --0150
  X"50", X"45", X"D2", X"46", X"4C", X"41", X"53", X"C8", --0158
  X"42", X"52", X"49", X"47", X"48", X"D4", X"49", X"4E", --0160
  X"56", X"45", X"52", X"53", X"C5", X"4F", X"56", X"45", --0168
  X"D2", X"4F", X"55", X"D4", X"4C", X"50", X"52", X"49", --0170
  X"4E", X"D4", X"4C", X"4C", X"49", X"53", X"D4", X"53", --0178
  X"54", X"4F", X"D0", X"52", X"45", X"41", X"C4", X"44", --0180
  X"41", X"54", X"C1", X"52", X"45", X"53", X"54", X"4F", --0188
  X"52", X"C5", X"4E", X"45", X"D7", X"42", X"4F", X"52", --0190
  X"44", X"45", X"D2", X"43", X"4F", X"4E", X"54", X"49", --0198
  X"4E", X"55", X"C5", X"44", X"49", X"CD", X"52", X"45", --01A0
  X"CD", X"46", X"4F", X"D2", X"47", X"4F", X"20", X"54", --01A8
  X"CF", X"47", X"4F", X"20", X"53", X"55", X"C2", X"49", --01B0
  X"4E", X"50", X"55", X"D4", X"4C", X"4F", X"41", X"C4", --01B8
  X"4C", X"49", X"53", X"D4", X"4C", X"45", X"D4", X"50", --01C0
  X"41", X"55", X"53", X"C5", X"4E", X"45", X"58", X"D4", --01C8
  X"50", X"4F", X"4B", X"C5", X"50", X"52", X"49", X"4E", --01D0
  X"D4", X"50", X"4C", X"4F", X"D4", X"52", X"55", X"CE", --01D8
  X"53", X"41", X"56", X"C5", X"52", X"41", X"4E", X"44", --01E0
  X"4F", X"4D", X"49", X"5A", X"C5", X"49", X"C6", X"43", --01E8
  X"4C", X"D3", X"44", X"52", X"41", X"D7", X"43", X"4C", --01F0
  X"45", X"41", X"D2", X"52", X"45", X"54", X"55", X"52", --01F8
  X"CE", X"43", X"4F", X"50", X"D9", X"42", X"48", X"59", --0200
  X"36", X"35", X"54", X"47", X"56", X"4E", X"4A", X"55", --0208
  X"37", X"34", X"52", X"46", X"43", X"4D", X"4B", X"49", --0210
  X"38", X"33", X"45", X"44", X"58", X"0E", X"4C", X"4F", --0218
  X"39", X"32", X"57", X"53", X"5A", X"20", X"0D", X"50", --0220
  X"30", X"31", X"51", X"41", X"E3", X"C4", X"E0", X"E4", --0228
  X"B4", X"BC", X"BD", X"BB", X"AF", X"B0", X"B1", X"C0", --0230
  X"A7", X"A6", X"BE", X"AD", X"B2", X"BA", X"E5", X"A5", --0238
  X"C2", X"E1", X"B3", X"B9", X"C1", X"B8", X"7E", X"DC", --0240
  X"DA", X"5C", X"B7", X"7B", X"7D", X"D8", X"BF", X"AE", --0248
  X"AA", X"AB", X"DD", X"DE", X"DF", X"7F", X"B5", X"D6", --0250
  X"7C", X"D5", X"5D", X"DB", X"B6", X"D9", X"5B", X"D7", --0258
  X"0C", X"07", X"06", X"04", X"05", X"08", X"0A", X"0B", --0260
  X"09", X"0F", X"E2", X"2A", X"3F", X"CD", X"C8", X"CC", --0268
  X"CB", X"5E", X"AC", X"2D", X"2B", X"3D", X"2E", X"2C", --0270
  X"3B", X"22", X"C7", X"3C", X"C3", X"3E", X"C5", X"2F", --0278
  X"C9", X"60", X"C6", X"3A", X"D0", X"CE", X"A8", X"CA", --0280
  X"D3", X"D4", X"D1", X"D2", X"A9", X"CF", X"2E", X"2F", --0288
  X"11", X"FF", X"FF", X"01", X"FE", X"FE", X"ED", X"78", --0290
  X"2F", X"E6", X"1F", X"28", X"0E", X"67", X"7D", X"14", --0298
  X"C0", X"D6", X"08", X"CB", X"3C", X"30", X"FA", X"53", --02A0
  X"5F", X"20", X"F4", X"2D", X"CB", X"00", X"38", X"E6", --02A8
  X"7A", X"3C", X"C8", X"FE", X"28", X"C8", X"FE", X"19", --02B0
  X"C8", X"7B", X"5A", X"57", X"FE", X"18", X"C9", X"CD", --02B8
  X"8E", X"02", X"C0", X"21", X"00", X"5C", X"CB", X"7E", --02C0
  X"20", X"07", X"23", X"35", X"2B", X"20", X"02", X"36", --02C8
  X"FF", X"7D", X"21", X"04", X"5C", X"BD", X"20", X"EE", --02D0
  X"CD", X"1E", X"03", X"D0", X"21", X"00", X"5C", X"BE", --02D8
  X"28", X"2E", X"EB", X"21", X"04", X"5C", X"BE", X"28", --02E0
  X"27", X"CB", X"7E", X"20", X"04", X"EB", X"CB", X"7E", --02E8
  X"C8", X"5F", X"77", X"23", X"36", X"05", X"23", X"3A", --02F0
  X"09", X"5C", X"77", X"23", X"FD", X"4E", X"07", X"FD", --02F8
  X"56", X"01", X"E5", X"CD", X"33", X"03", X"E1", X"77", --0300
  X"32", X"08", X"5C", X"FD", X"CB", X"01", X"EE", X"C9", --0308
  X"23", X"36", X"05", X"23", X"35", X"C0", X"3A", X"0A", --0310
  X"5C", X"77", X"23", X"7E", X"18", X"EA", X"42", X"16", --0318
  X"00", X"7B", X"FE", X"27", X"D0", X"FE", X"18", X"20", --0320
  X"03", X"CB", X"78", X"C0", X"21", X"05", X"02", X"19", --0328
  X"7E", X"37", X"C9", X"7B", X"FE", X"3A", X"38", X"2F", --0330
  X"0D", X"FA", X"4F", X"03", X"28", X"03", X"C6", X"4F", --0338
  X"C9", X"21", X"EB", X"01", X"04", X"28", X"03", X"21", --0340
  X"05", X"02", X"16", X"00", X"19", X"7E", X"C9", X"21", --0348
  X"29", X"02", X"CB", X"40", X"28", X"F4", X"CB", X"5A", --0350
  X"28", X"0A", X"FD", X"CB", X"30", X"5E", X"C0", X"04", --0358
  X"C0", X"C6", X"20", X"C9", X"C6", X"A5", X"C9", X"FE", --0360
  X"30", X"D8", X"0D", X"FA", X"9D", X"03", X"20", X"19", --0368
  X"21", X"54", X"02", X"CB", X"68", X"28", X"D3", X"FE", --0370
  X"38", X"30", X"07", X"D6", X"20", X"04", X"C8", X"C6", --0378
  X"08", X"C9", X"D6", X"36", X"04", X"C8", X"C6", X"FE", --0380
  X"C9", X"21", X"30", X"02", X"FE", X"39", X"28", X"BA", --0388
  X"FE", X"30", X"28", X"B6", X"E6", X"07", X"C6", X"80", --0390
  X"04", X"C8", X"EE", X"0F", X"C9", X"04", X"C8", X"CB", --0398
  X"68", X"21", X"30", X"02", X"20", X"A4", X"D6", X"10", --03A0
  X"FE", X"22", X"28", X"06", X"FE", X"20", X"C0", X"3E", --03A8
  X"5F", X"C9", X"3E", X"40", X"C9", X"F3", X"7D", X"CB", --03B0
  X"3D", X"CB", X"3D", X"2F", X"E6", X"03", X"4F", X"06", --03B8
  X"00", X"DD", X"21", X"D1", X"03", X"DD", X"09", X"3A", --03C0
  X"48", X"5C", X"E6", X"38", X"0F", X"0F", X"0F", X"F6", --03C8
  X"08", X"00", X"00", X"00", X"04", X"0C", X"0D", X"20", --03D0
  X"FD", X"0E", X"3F", X"05", X"C2", X"D6", X"03", X"EE", --03D8
  X"10", X"D3", X"FE", X"44", X"4F", X"CB", X"67", X"20", --03E0
  X"09", X"7A", X"B3", X"28", X"09", X"79", X"4D", X"1B", --03E8
  X"DD", X"E9", X"4D", X"0C", X"DD", X"E9", X"FB", X"C9", --03F0
  X"EF", X"31", X"27", X"C0", X"03", X"34", X"EC", X"6C", --03F8
  X"98", X"1F", X"F5", X"04", X"A1", X"0F", X"38", X"21", --0400
  X"92", X"5C", X"7E", X"A7", X"20", X"5E", X"23", X"4E", --0408
  X"23", X"46", X"78", X"17", X"9F", X"B9", X"20", X"54", --0410
  X"23", X"BE", X"20", X"50", X"78", X"C6", X"3C", X"F2", --0418
  X"25", X"04", X"E2", X"6C", X"04", X"06", X"FA", X"04", --0420
  X"D6", X"0C", X"30", X"FB", X"C6", X"0C", X"C5", X"21", --0428
  X"6E", X"04", X"CD", X"06", X"34", X"CD", X"B4", X"33", --0430
  X"EF", X"04", X"38", X"F1", X"86", X"77", X"EF", X"C0", --0438
  X"02", X"31", X"38", X"CD", X"94", X"1E", X"FE", X"0B", --0440
  X"30", X"22", X"EF", X"E0", X"04", X"E0", X"34", X"80", --0448
  X"43", X"55", X"9F", X"80", X"01", X"05", X"34", X"35", --0450
  X"71", X"03", X"38", X"CD", X"99", X"1E", X"C5", X"CD", --0458
  X"99", X"1E", X"E1", X"50", X"59", X"7A", X"B3", X"C8", --0460
  X"1B", X"C3", X"B5", X"03", X"CF", X"0A", X"89", X"02", --0468
  X"D0", X"12", X"86", X"89", X"0A", X"97", X"60", X"75", --0470
  X"89", X"12", X"D5", X"17", X"1F", X"89", X"1B", X"90", --0478
  X"41", X"02", X"89", X"24", X"D0", X"53", X"CA", X"89", --0480
  X"2E", X"9D", X"36", X"B1", X"89", X"38", X"FF", X"49", --0488
  X"3E", X"89", X"43", X"FF", X"6A", X"73", X"89", X"4F", --0490
  X"A7", X"00", X"54", X"89", X"5C", X"00", X"00", X"00", --0498
  X"89", X"69", X"14", X"F6", X"24", X"89", X"76", X"F1", --04A0
  X"10", X"05", X"CD", X"FB", X"24", X"3A", X"3B", X"5C", --04A8
  X"87", X"FA", X"8A", X"1C", X"E1", X"D0", X"E5", X"CD", --04B0
  X"F1", X"2B", X"62", X"6B", X"0D", X"F8", X"09", X"CB", --04B8
  X"FE", X"C9", X"21", X"3F", X"05", X"E5", X"21", X"80", --04C0
  X"1F", X"CB", X"7F", X"28", X"03", X"21", X"98", X"0C", --04C8
  X"08", X"13", X"DD", X"2B", X"F3", X"3E", X"02", X"47", --04D0
  X"10", X"FE", X"D3", X"FE", X"EE", X"0F", X"06", X"A4", --04D8
  X"2D", X"20", X"F5", X"05", X"25", X"F2", X"D8", X"04", --04E0
  X"06", X"2F", X"10", X"FE", X"D3", X"FE", X"3E", X"0D", --04E8
  X"06", X"37", X"10", X"FE", X"D3", X"FE", X"01", X"0E", --04F0
  X"3B", X"08", X"6F", X"C3", X"07", X"05", X"7A", X"B3", --04F8
  X"28", X"0C", X"DD", X"6E", X"00", X"7C", X"AD", X"67", --0500
  X"3E", X"01", X"37", X"C3", X"25", X"05", X"6C", X"18", --0508
  X"F4", X"79", X"CB", X"78", X"10", X"FE", X"30", X"04", --0510
  X"06", X"42", X"10", X"FE", X"D3", X"FE", X"06", X"3E", --0518
  X"20", X"EF", X"05", X"AF", X"3C", X"CB", X"15", X"C2", --0520
  X"14", X"05", X"1B", X"DD", X"23", X"06", X"31", X"3E", --0528
  X"7F", X"DB", X"FE", X"1F", X"D0", X"7A", X"3C", X"C2", --0530
  X"FE", X"04", X"06", X"3B", X"10", X"FE", X"C9", X"F5", --0538
  X"3A", X"48", X"5C", X"E6", X"38", X"0F", X"0F", X"0F", --0540
  X"D3", X"FE", X"3E", X"7F", X"DB", X"FE", X"1F", X"FB", --0548
  X"38", X"02", X"CF", X"0C", X"F1", X"C9", X"14", X"08", --0550
  X"15", X"F3", X"3E", X"0F", X"D3", X"FE", X"21", X"3F", --0558
  X"05", X"E5", X"DB", X"FE", X"1F", X"E6", X"20", X"F6", --0560
  X"02", X"4F", X"BF", X"C0", X"CD", X"E7", X"05", X"30", --0568
  X"FA", X"21", X"15", X"04", X"10", X"FE", X"2B", X"7C", --0570
  X"B5", X"20", X"F9", X"CD", X"E3", X"05", X"30", X"EB", --0578
  X"06", X"9C", X"CD", X"E3", X"05", X"30", X"E4", X"3E", --0580
  X"C6", X"B8", X"30", X"E0", X"24", X"20", X"F1", X"06", --0588
  X"C9", X"CD", X"E7", X"05", X"30", X"D5", X"78", X"FE", --0590
  X"D4", X"30", X"F4", X"CD", X"E7", X"05", X"D0", X"79", --0598
  X"EE", X"03", X"4F", X"26", X"00", X"06", X"B0", X"18", --05A0
  X"1F", X"08", X"20", X"07", X"30", X"0F", X"DD", X"75", --05A8
  X"00", X"18", X"0F", X"CB", X"11", X"AD", X"C0", X"79", --05B0
  X"1F", X"4F", X"13", X"18", X"07", X"DD", X"7E", X"00", --05B8
  X"AD", X"C0", X"DD", X"23", X"1B", X"08", X"06", X"B2", --05C0
  X"2E", X"01", X"CD", X"E3", X"05", X"D0", X"3E", X"CB", --05C8
  X"B8", X"CB", X"15", X"06", X"B0", X"D2", X"CA", X"05", --05D0
  X"7C", X"AD", X"67", X"7A", X"B3", X"20", X"CA", X"7C", --05D8
  X"FE", X"01", X"C9", X"CD", X"E7", X"05", X"D0", X"3E", --05E0
  X"16", X"3D", X"20", X"FD", X"A7", X"04", X"C8", X"3E", --05E8
  X"7F", X"DB", X"FE", X"1F", X"D0", X"A9", X"E6", X"20", --05F0
  X"28", X"F3", X"79", X"2F", X"4F", X"E6", X"07", X"F6", --05F8
  X"08", X"D3", X"FE", X"37", X"C9", X"F1", X"3A", X"74", --0600
  X"5C", X"D6", X"E0", X"32", X"74", X"5C", X"CD", X"8C", --0608
  X"1C", X"CD", X"30", X"25", X"28", X"3C", X"01", X"11", --0610
  X"00", X"3A", X"74", X"5C", X"A7", X"28", X"02", X"0E", --0618
  X"22", X"F7", X"D5", X"DD", X"E1", X"06", X"0B", X"3E", --0620
  X"20", X"12", X"13", X"10", X"FC", X"DD", X"36", X"01", --0628
  X"FF", X"CD", X"F1", X"2B", X"21", X"F6", X"FF", X"0B", --0630
  X"09", X"03", X"30", X"0F", X"3A", X"74", X"5C", X"A7", --0638
  X"20", X"02", X"CF", X"0E", X"78", X"B1", X"28", X"0A", --0640
  X"01", X"0A", X"00", X"DD", X"E5", X"E1", X"23", X"EB", --0648
  X"ED", X"B0", X"DF", X"FE", X"E4", X"20", X"49", X"3A", --0650
  X"74", X"5C", X"FE", X"03", X"CA", X"8A", X"1C", X"E7", --0658
  X"CD", X"B2", X"28", X"CB", X"F9", X"30", X"0B", X"21", --0660
  X"00", X"00", X"3A", X"74", X"5C", X"3D", X"28", X"15", --0668
  X"CF", X"01", X"C2", X"8A", X"1C", X"CD", X"30", X"25", --0670
  X"28", X"18", X"23", X"7E", X"DD", X"77", X"0B", X"23", --0678
  X"7E", X"DD", X"77", X"0C", X"23", X"DD", X"71", X"0E", --0680
  X"3E", X"01", X"CB", X"71", X"28", X"01", X"3C", X"DD", --0688
  X"77", X"00", X"EB", X"E7", X"FE", X"29", X"20", X"DA", --0690
  X"E7", X"CD", X"EE", X"1B", X"EB", X"C3", X"5A", X"07", --0698
  X"FE", X"AA", X"20", X"1F", X"3A", X"74", X"5C", X"FE", --06A0
  X"03", X"CA", X"8A", X"1C", X"E7", X"CD", X"EE", X"1B", --06A8
  X"DD", X"36", X"0B", X"00", X"DD", X"36", X"0C", X"1B", --06B0
  X"21", X"00", X"40", X"DD", X"75", X"0D", X"DD", X"74", --06B8
  X"0E", X"18", X"4D", X"FE", X"AF", X"20", X"4F", X"3A", --06C0
  X"74", X"5C", X"FE", X"03", X"CA", X"8A", X"1C", X"E7", --06C8
  X"CD", X"48", X"20", X"20", X"0C", X"3A", X"74", X"5C", --06D0
  X"A7", X"CA", X"8A", X"1C", X"CD", X"E6", X"1C", X"18", --06D8
  X"0F", X"CD", X"82", X"1C", X"DF", X"FE", X"2C", X"28", --06E0
  X"0C", X"3A", X"74", X"5C", X"A7", X"CA", X"8A", X"1C", --06E8
  X"CD", X"E6", X"1C", X"18", X"04", X"E7", X"CD", X"82", --06F0
  X"1C", X"CD", X"EE", X"1B", X"CD", X"99", X"1E", X"DD", --06F8
  X"71", X"0B", X"DD", X"70", X"0C", X"CD", X"99", X"1E", --0700
  X"DD", X"71", X"0D", X"DD", X"70", X"0E", X"60", X"69", --0708
  X"DD", X"36", X"00", X"03", X"18", X"44", X"FE", X"CA", --0710
  X"28", X"09", X"CD", X"EE", X"1B", X"DD", X"36", X"0E", --0718
  X"80", X"18", X"17", X"3A", X"74", X"5C", X"A7", X"C2", --0720
  X"8A", X"1C", X"E7", X"CD", X"82", X"1C", X"CD", X"EE", --0728
  X"1B", X"CD", X"99", X"1E", X"DD", X"71", X"0D", X"DD", --0730
  X"70", X"0E", X"DD", X"36", X"00", X"00", X"2A", X"59", --0738
  X"5C", X"ED", X"5B", X"53", X"5C", X"37", X"ED", X"52", --0740
  X"DD", X"75", X"0B", X"DD", X"74", X"0C", X"2A", X"4B", --0748
  X"5C", X"ED", X"52", X"DD", X"75", X"0F", X"DD", X"74", --0750
  X"10", X"EB", X"3A", X"74", X"5C", X"A7", X"CA", X"70", --0758
  X"09", X"E5", X"01", X"11", X"00", X"DD", X"09", X"DD", --0760
  X"E5", X"11", X"11", X"00", X"AF", X"37", X"CD", X"56", --0768
  X"05", X"DD", X"E1", X"30", X"F2", X"3E", X"FE", X"CD", --0770
  X"01", X"16", X"FD", X"36", X"52", X"03", X"0E", X"80", --0778
  X"DD", X"7E", X"00", X"DD", X"BE", X"EF", X"20", X"02", --0780
  X"0E", X"F6", X"FE", X"04", X"30", X"D9", X"11", X"C0", --0788
  X"09", X"C5", X"CD", X"0A", X"0C", X"C1", X"DD", X"E5", --0790
  X"D1", X"21", X"F0", X"FF", X"19", X"06", X"0A", X"7E", --0798
  X"3C", X"20", X"03", X"79", X"80", X"4F", X"13", X"1A", --07A0
  X"BE", X"23", X"20", X"01", X"0C", X"D7", X"10", X"F6", --07A8
  X"CB", X"79", X"20", X"B3", X"3E", X"0D", X"D7", X"E1", --07B0
  X"DD", X"7E", X"00", X"FE", X"03", X"28", X"0C", X"3A", --07B8
  X"74", X"5C", X"3D", X"CA", X"08", X"08", X"FE", X"02", --07C0
  X"CA", X"B6", X"08", X"E5", X"DD", X"6E", X"FA", X"DD", --07C8
  X"66", X"FB", X"DD", X"5E", X"0B", X"DD", X"56", X"0C", --07D0
  X"7C", X"B5", X"28", X"0D", X"ED", X"52", X"38", X"26", --07D8
  X"28", X"07", X"DD", X"7E", X"00", X"FE", X"03", X"20", --07E0
  X"1D", X"E1", X"7C", X"B5", X"20", X"06", X"DD", X"6E", --07E8
  X"0D", X"DD", X"66", X"0E", X"E5", X"DD", X"E1", X"3A", --07F0
  X"74", X"5C", X"FE", X"02", X"37", X"20", X"01", X"A7", --07F8
  X"3E", X"FF", X"CD", X"56", X"05", X"D8", X"CF", X"1A", --0800
  X"DD", X"5E", X"0B", X"DD", X"56", X"0C", X"E5", X"7C", --0808
  X"B5", X"20", X"06", X"13", X"13", X"13", X"EB", X"18", --0810
  X"0C", X"DD", X"6E", X"FA", X"DD", X"66", X"FB", X"EB", --0818
  X"37", X"ED", X"52", X"38", X"09", X"11", X"05", X"00", --0820
  X"19", X"44", X"4D", X"CD", X"05", X"1F", X"E1", X"DD", --0828
  X"7E", X"00", X"A7", X"28", X"3E", X"7C", X"B5", X"28", --0830
  X"13", X"2B", X"46", X"2B", X"4E", X"2B", X"03", X"03", --0838
  X"03", X"DD", X"22", X"5F", X"5C", X"CD", X"E8", X"19", --0840
  X"DD", X"2A", X"5F", X"5C", X"2A", X"59", X"5C", X"2B", --0848
  X"DD", X"4E", X"0B", X"DD", X"46", X"0C", X"C5", X"03", --0850
  X"03", X"03", X"DD", X"7E", X"FD", X"F5", X"CD", X"55", --0858
  X"16", X"23", X"F1", X"77", X"D1", X"23", X"73", X"23", --0860
  X"72", X"23", X"E5", X"DD", X"E1", X"37", X"3E", X"FF", --0868
  X"C3", X"02", X"08", X"EB", X"2A", X"59", X"5C", X"2B", --0870
  X"DD", X"22", X"5F", X"5C", X"DD", X"4E", X"0B", X"DD", --0878
  X"46", X"0C", X"C5", X"CD", X"E5", X"19", X"C1", X"E5", --0880
  X"C5", X"CD", X"55", X"16", X"DD", X"2A", X"5F", X"5C", --0888
  X"23", X"DD", X"4E", X"0F", X"DD", X"46", X"10", X"09", --0890
  X"22", X"4B", X"5C", X"DD", X"66", X"0E", X"7C", X"E6", --0898
  X"C0", X"20", X"0A", X"DD", X"6E", X"0D", X"22", X"42", --08A0
  X"5C", X"FD", X"36", X"0A", X"00", X"D1", X"DD", X"E1", --08A8
  X"37", X"3E", X"FF", X"C3", X"02", X"08", X"DD", X"4E", --08B0
  X"0B", X"DD", X"46", X"0C", X"C5", X"03", X"F7", X"36", --08B8
  X"80", X"EB", X"D1", X"E5", X"E5", X"DD", X"E1", X"37", --08C0
  X"3E", X"FF", X"CD", X"02", X"08", X"E1", X"ED", X"5B", --08C8
  X"53", X"5C", X"7E", X"E6", X"C0", X"20", X"19", X"1A", --08D0
  X"13", X"BE", X"23", X"20", X"02", X"1A", X"BE", X"1B", --08D8
  X"2B", X"30", X"08", X"E5", X"EB", X"CD", X"B8", X"19", --08E0
  X"E1", X"18", X"EC", X"CD", X"2C", X"09", X"18", X"E2", --08E8
  X"7E", X"4F", X"FE", X"80", X"C8", X"E5", X"2A", X"4B", --08F0
  X"5C", X"7E", X"FE", X"80", X"28", X"25", X"B9", X"28", --08F8
  X"08", X"C5", X"CD", X"B8", X"19", X"C1", X"EB", X"18", --0900
  X"F0", X"E6", X"E0", X"FE", X"A0", X"20", X"12", X"D1", --0908
  X"D5", X"E5", X"23", X"13", X"1A", X"BE", X"20", X"06", --0910
  X"17", X"30", X"F7", X"E1", X"18", X"03", X"E1", X"18", --0918
  X"E0", X"3E", X"FF", X"D1", X"EB", X"3C", X"37", X"CD", --0920
  X"2C", X"09", X"18", X"C4", X"20", X"10", X"08", X"22", --0928
  X"5F", X"5C", X"EB", X"CD", X"B8", X"19", X"CD", X"E8", --0930
  X"19", X"EB", X"2A", X"5F", X"5C", X"08", X"08", X"D5", --0938
  X"CD", X"B8", X"19", X"22", X"5F", X"5C", X"2A", X"53", --0940
  X"5C", X"E3", X"C5", X"08", X"38", X"07", X"2B", X"CD", --0948
  X"55", X"16", X"23", X"18", X"03", X"CD", X"55", X"16", --0950
  X"23", X"C1", X"D1", X"ED", X"53", X"53", X"5C", X"ED", --0958
  X"5B", X"5F", X"5C", X"C5", X"D5", X"EB", X"ED", X"B0", --0960
  X"E1", X"C1", X"D5", X"CD", X"E8", X"19", X"D1", X"C9", --0968
  X"E5", X"3E", X"FD", X"CD", X"01", X"16", X"AF", X"11", --0970
  X"A1", X"09", X"CD", X"0A", X"0C", X"FD", X"CB", X"02", --0978
  X"EE", X"CD", X"D4", X"15", X"DD", X"E5", X"11", X"11", --0980
  X"00", X"AF", X"CD", X"C2", X"04", X"DD", X"E1", X"06", --0988
  X"32", X"76", X"10", X"FD", X"DD", X"5E", X"0B", X"DD", --0990
  X"56", X"0C", X"3E", X"FF", X"DD", X"E1", X"C3", X"C2", --0998
  X"04", X"80", X"53", X"74", X"61", X"72", X"74", X"20", --09A0
  X"74", X"61", X"70", X"65", X"2C", X"20", X"74", X"68", --09A8
  X"65", X"6E", X"20", X"70", X"72", X"65", X"73", X"73", --09B0
  X"20", X"61", X"6E", X"79", X"20", X"6B", X"65", X"79", --09B8
  X"AE", X"0D", X"50", X"72", X"6F", X"67", X"72", X"61", --09C0
  X"6D", X"3A", X"A0", X"0D", X"4E", X"75", X"6D", X"62", --09C8
  X"65", X"72", X"20", X"61", X"72", X"72", X"61", X"79", --09D0
  X"3A", X"A0", X"0D", X"43", X"68", X"61", X"72", X"61", --09D8
  X"63", X"74", X"65", X"72", X"20", X"61", X"72", X"72", --09E0
  X"61", X"79", X"3A", X"A0", X"0D", X"42", X"79", X"74", --09E8
  X"65", X"73", X"3A", X"A0", X"CD", X"03", X"0B", X"FE", --09F0
  X"20", X"D2", X"D9", X"0A", X"FE", X"06", X"38", X"69", --09F8
  X"FE", X"18", X"30", X"65", X"21", X"0B", X"0A", X"5F", --0A00
  X"16", X"00", X"19", X"5E", X"19", X"E5", X"C3", X"03", --0A08
  X"0B", X"4E", X"57", X"10", X"29", X"54", X"53", X"52", --0A10
  X"37", X"50", X"4F", X"5F", X"5E", X"5D", X"5C", X"5B", --0A18
  X"5A", X"54", X"53", X"0C", X"3E", X"22", X"B9", X"20", --0A20
  X"11", X"FD", X"CB", X"01", X"4E", X"20", X"09", X"04", --0A28
  X"0E", X"02", X"3E", X"18", X"B8", X"20", X"03", X"05", --0A30
  X"0E", X"21", X"C3", X"D9", X"0D", X"3A", X"91", X"5C", --0A38
  X"F5", X"FD", X"36", X"57", X"01", X"3E", X"20", X"CD", --0A40
  X"65", X"0B", X"F1", X"32", X"91", X"5C", X"C9", X"FD", --0A48
  X"CB", X"01", X"4E", X"C2", X"CD", X"0E", X"0E", X"21", --0A50
  X"CD", X"55", X"0C", X"05", X"C3", X"D9", X"0D", X"CD", --0A58
  X"03", X"0B", X"79", X"3D", X"3D", X"E6", X"10", X"18", --0A60
  X"5A", X"3E", X"3F", X"18", X"6C", X"11", X"87", X"0A", --0A68
  X"32", X"0F", X"5C", X"18", X"0B", X"11", X"6D", X"0A", --0A70
  X"18", X"03", X"11", X"87", X"0A", X"32", X"0E", X"5C", --0A78
  X"2A", X"51", X"5C", X"73", X"23", X"72", X"C9", X"11", --0A80
  X"F4", X"09", X"CD", X"80", X"0A", X"2A", X"0E", X"5C", --0A88
  X"57", X"7D", X"FE", X"16", X"DA", X"11", X"22", X"20", --0A90
  X"29", X"44", X"4A", X"3E", X"1F", X"91", X"38", X"0C", --0A98
  X"C6", X"02", X"4F", X"FD", X"CB", X"01", X"4E", X"20", --0AA0
  X"16", X"3E", X"16", X"90", X"DA", X"9F", X"1E", X"3C", --0AA8
  X"47", X"04", X"FD", X"CB", X"02", X"46", X"C2", X"55", --0AB0
  X"0C", X"FD", X"BE", X"31", X"DA", X"86", X"0C", X"C3", --0AB8
  X"D9", X"0D", X"7C", X"CD", X"03", X"0B", X"81", X"3D", --0AC0
  X"E6", X"1F", X"C8", X"57", X"FD", X"CB", X"01", X"C6", --0AC8
  X"3E", X"20", X"CD", X"3B", X"0C", X"15", X"20", X"F8", --0AD0
  X"C9", X"CD", X"24", X"0B", X"FD", X"CB", X"01", X"4E", --0AD8
  X"20", X"1A", X"FD", X"CB", X"02", X"46", X"20", X"08", --0AE0
  X"ED", X"43", X"88", X"5C", X"22", X"84", X"5C", X"C9", --0AE8
  X"ED", X"43", X"8A", X"5C", X"ED", X"43", X"82", X"5C", --0AF0
  X"22", X"86", X"5C", X"C9", X"FD", X"71", X"45", X"22", --0AF8
  X"80", X"5C", X"C9", X"FD", X"CB", X"01", X"4E", X"20", --0B00
  X"14", X"ED", X"4B", X"88", X"5C", X"2A", X"84", X"5C", --0B08
  X"FD", X"CB", X"02", X"46", X"C8", X"ED", X"4B", X"8A", --0B10
  X"5C", X"2A", X"86", X"5C", X"C9", X"FD", X"4E", X"45", --0B18
  X"2A", X"80", X"5C", X"C9", X"FE", X"80", X"38", X"3D", --0B20
  X"FE", X"90", X"30", X"26", X"47", X"CD", X"38", X"0B", --0B28
  X"CD", X"03", X"0B", X"11", X"92", X"5C", X"18", X"47", --0B30
  X"21", X"92", X"5C", X"CD", X"3E", X"0B", X"CB", X"18", --0B38
  X"9F", X"E6", X"0F", X"4F", X"CB", X"18", X"9F", X"E6", --0B40
  X"F0", X"B1", X"0E", X"04", X"77", X"23", X"0D", X"20", --0B48
  X"FB", X"C9", X"D6", X"A5", X"30", X"09", X"C6", X"15", --0B50
  X"C5", X"ED", X"4B", X"7B", X"5C", X"18", X"0B", X"CD", --0B58
  X"10", X"0C", X"C3", X"03", X"0B", X"C5", X"ED", X"4B", --0B60
  X"36", X"5C", X"EB", X"21", X"3B", X"5C", X"CB", X"86", --0B68
  X"FE", X"20", X"20", X"02", X"CB", X"C6", X"26", X"00", --0B70
  X"6F", X"29", X"29", X"29", X"09", X"C1", X"EB", X"79", --0B78
  X"3D", X"3E", X"21", X"20", X"0E", X"05", X"4F", X"FD", --0B80
  X"CB", X"01", X"4E", X"28", X"06", X"D5", X"CD", X"CD", --0B88
  X"0E", X"D1", X"79", X"B9", X"D5", X"CC", X"55", X"0C", --0B90
  X"D1", X"C5", X"E5", X"3A", X"91", X"5C", X"06", X"FF", --0B98
  X"1F", X"38", X"01", X"04", X"1F", X"1F", X"9F", X"4F", --0BA0
  X"3E", X"08", X"A7", X"FD", X"CB", X"01", X"4E", X"28", --0BA8
  X"05", X"FD", X"CB", X"30", X"CE", X"37", X"EB", X"08", --0BB0
  X"1A", X"A0", X"AE", X"A9", X"12", X"08", X"38", X"13", --0BB8
  X"14", X"23", X"3D", X"20", X"F2", X"EB", X"25", X"FD", --0BC0
  X"CB", X"01", X"4E", X"CC", X"DB", X"0B", X"E1", X"C1", --0BC8
  X"0D", X"23", X"C9", X"08", X"3E", X"20", X"83", X"5F", --0BD0
  X"08", X"18", X"E6", X"7C", X"0F", X"0F", X"0F", X"E6", --0BD8
  X"03", X"F6", X"58", X"67", X"ED", X"5B", X"8F", X"5C", --0BE0
  X"7E", X"AB", X"A2", X"AB", X"FD", X"CB", X"57", X"76", --0BE8
  X"28", X"08", X"E6", X"C7", X"CB", X"57", X"20", X"02", --0BF0
  X"EE", X"38", X"FD", X"CB", X"57", X"66", X"28", X"08", --0BF8
  X"E6", X"F8", X"CB", X"6F", X"20", X"02", X"EE", X"07", --0C00
  X"77", X"C9", X"E5", X"26", X"00", X"E3", X"18", X"04", --0C08
  X"11", X"95", X"00", X"F5", X"CD", X"41", X"0C", X"38", --0C10
  X"09", X"3E", X"20", X"FD", X"CB", X"01", X"46", X"CC", --0C18
  X"3B", X"0C", X"1A", X"E6", X"7F", X"CD", X"3B", X"0C", --0C20
  X"1A", X"13", X"87", X"30", X"F5", X"D1", X"FE", X"48", --0C28
  X"28", X"03", X"FE", X"82", X"D8", X"7A", X"FE", X"03", --0C30
  X"D8", X"3E", X"20", X"D5", X"D9", X"D7", X"D9", X"D1", --0C38
  X"C9", X"F5", X"EB", X"3C", X"CB", X"7E", X"23", X"28", --0C40
  X"FB", X"3D", X"20", X"F8", X"EB", X"F1", X"FE", X"20", --0C48
  X"D8", X"1A", X"D6", X"41", X"C9", X"FD", X"CB", X"01", --0C50
  X"4E", X"C0", X"11", X"D9", X"0D", X"D5", X"78", X"FD", --0C58
  X"CB", X"02", X"46", X"C2", X"02", X"0D", X"FD", X"BE", --0C60
  X"31", X"38", X"1B", X"C0", X"FD", X"CB", X"02", X"66", --0C68
  X"28", X"16", X"FD", X"5E", X"2D", X"1D", X"28", X"5A", --0C70
  X"3E", X"00", X"CD", X"01", X"16", X"ED", X"7B", X"3F", --0C78
  X"5C", X"FD", X"CB", X"02", X"A6", X"C9", X"CF", X"04", --0C80
  X"FD", X"35", X"52", X"20", X"45", X"3E", X"18", X"90", --0C88
  X"32", X"8C", X"5C", X"2A", X"8F", X"5C", X"E5", X"3A", --0C90
  X"91", X"5C", X"F5", X"3E", X"FD", X"CD", X"01", X"16", --0C98
  X"AF", X"11", X"F8", X"0C", X"CD", X"0A", X"0C", X"FD", --0CA0
  X"CB", X"02", X"EE", X"21", X"3B", X"5C", X"CB", X"DE", --0CA8
  X"CB", X"AE", X"D9", X"CD", X"D4", X"15", X"D9", X"FE", --0CB0
  X"20", X"28", X"45", X"FE", X"E2", X"28", X"41", X"F6", --0CB8
  X"20", X"FE", X"6E", X"28", X"3B", X"3E", X"FE", X"CD", --0CC0
  X"01", X"16", X"F1", X"32", X"91", X"5C", X"E1", X"22", --0CC8
  X"8F", X"5C", X"CD", X"FE", X"0D", X"FD", X"46", X"31", --0CD0
  X"04", X"0E", X"21", X"C5", X"CD", X"9B", X"0E", X"7C", --0CD8
  X"0F", X"0F", X"0F", X"E6", X"03", X"F6", X"58", X"67", --0CE0
  X"11", X"E0", X"5A", X"1A", X"4E", X"06", X"20", X"EB", --0CE8
  X"12", X"71", X"13", X"23", X"10", X"FA", X"C1", X"C9", --0CF0
  X"80", X"73", X"63", X"72", X"6F", X"6C", X"6C", X"BF", --0CF8
  X"CF", X"0C", X"FE", X"02", X"38", X"80", X"FD", X"86", --0D00
  X"31", X"D6", X"19", X"D0", X"ED", X"44", X"C5", X"47", --0D08
  X"2A", X"8F", X"5C", X"E5", X"2A", X"91", X"5C", X"E5", --0D10
  X"CD", X"4D", X"0D", X"78", X"F5", X"21", X"6B", X"5C", --0D18
  X"46", X"78", X"3C", X"77", X"21", X"89", X"5C", X"BE", --0D20
  X"38", X"03", X"34", X"06", X"18", X"CD", X"00", X"0E", --0D28
  X"F1", X"3D", X"20", X"E8", X"E1", X"FD", X"75", X"57", --0D30
  X"E1", X"22", X"8F", X"5C", X"ED", X"4B", X"88", X"5C", --0D38
  X"FD", X"CB", X"02", X"86", X"CD", X"D9", X"0D", X"FD", --0D40
  X"CB", X"02", X"C6", X"C1", X"C9", X"AF", X"2A", X"8D", --0D48
  X"5C", X"FD", X"CB", X"02", X"46", X"28", X"04", X"67", --0D50
  X"FD", X"6E", X"0E", X"22", X"8F", X"5C", X"21", X"91", --0D58
  X"5C", X"20", X"02", X"7E", X"0F", X"AE", X"E6", X"55", --0D60
  X"AE", X"77", X"C9", X"CD", X"AF", X"0D", X"21", X"3C", --0D68
  X"5C", X"CB", X"AE", X"CB", X"C6", X"CD", X"4D", X"0D", --0D70
  X"FD", X"46", X"31", X"CD", X"44", X"0E", X"21", X"C0", --0D78
  X"5A", X"3A", X"8D", X"5C", X"05", X"18", X"07", X"0E", --0D80
  X"20", X"2B", X"77", X"0D", X"20", X"FB", X"10", X"F7", --0D88
  X"FD", X"36", X"31", X"02", X"3E", X"FD", X"CD", X"01", --0D90
  X"16", X"2A", X"51", X"5C", X"11", X"F4", X"09", X"A7", --0D98
  X"73", X"23", X"72", X"23", X"11", X"A8", X"10", X"3F", --0DA0
  X"38", X"F6", X"01", X"21", X"17", X"18", X"2A", X"21", --0DA8
  X"00", X"00", X"22", X"7D", X"5C", X"FD", X"CB", X"30", --0DB0
  X"86", X"CD", X"94", X"0D", X"3E", X"FE", X"CD", X"01", --0DB8
  X"16", X"CD", X"4D", X"0D", X"06", X"18", X"CD", X"44", --0DC0
  X"0E", X"2A", X"51", X"5C", X"11", X"F4", X"09", X"73", --0DC8
  X"23", X"72", X"FD", X"36", X"52", X"01", X"01", X"21", --0DD0
  X"18", X"21", X"00", X"5B", X"FD", X"CB", X"01", X"4E", --0DD8
  X"20", X"12", X"78", X"FD", X"CB", X"02", X"46", X"28", --0DE0
  X"05", X"FD", X"86", X"31", X"D6", X"18", X"C5", X"47", --0DE8
  X"CD", X"9B", X"0E", X"C1", X"3E", X"21", X"91", X"5F", --0DF0
  X"16", X"00", X"19", X"C3", X"DC", X"0A", X"06", X"17", --0DF8
  X"CD", X"9B", X"0E", X"0E", X"08", X"C5", X"E5", X"78", --0E00
  X"E6", X"07", X"78", X"20", X"0C", X"EB", X"21", X"E0", --0E08
  X"F8", X"19", X"EB", X"01", X"20", X"00", X"3D", X"ED", --0E10
  X"B0", X"EB", X"21", X"E0", X"FF", X"19", X"EB", X"47", --0E18
  X"E6", X"07", X"0F", X"0F", X"0F", X"4F", X"78", X"06", --0E20
  X"00", X"ED", X"B0", X"06", X"07", X"09", X"E6", X"F8", --0E28
  X"20", X"DB", X"E1", X"24", X"C1", X"0D", X"20", X"CD", --0E30
  X"CD", X"88", X"0E", X"21", X"E0", X"FF", X"19", X"EB", --0E38
  X"ED", X"B0", X"06", X"01", X"C5", X"CD", X"9B", X"0E", --0E40
  X"0E", X"08", X"C5", X"E5", X"78", X"E6", X"07", X"0F", --0E48
  X"0F", X"0F", X"4F", X"78", X"06", X"00", X"0D", X"54", --0E50
  X"5D", X"36", X"00", X"13", X"ED", X"B0", X"11", X"01", --0E58
  X"07", X"19", X"3D", X"E6", X"F8", X"47", X"20", X"E5", --0E60
  X"E1", X"24", X"C1", X"0D", X"20", X"DC", X"CD", X"88", --0E68
  X"0E", X"62", X"6B", X"13", X"3A", X"8D", X"5C", X"FD", --0E70
  X"CB", X"02", X"46", X"28", X"03", X"3A", X"48", X"5C", --0E78
  X"77", X"0B", X"ED", X"B0", X"C1", X"0E", X"21", X"C9", --0E80
  X"7C", X"0F", X"0F", X"0F", X"3D", X"F6", X"50", X"67", --0E88
  X"EB", X"61", X"68", X"29", X"29", X"29", X"29", X"29", --0E90
  X"44", X"4D", X"C9", X"3E", X"18", X"90", X"57", X"0F", --0E98
  X"0F", X"0F", X"E6", X"E0", X"6F", X"7A", X"E6", X"18", --0EA0
  X"F6", X"40", X"67", X"C9", X"F3", X"06", X"B0", X"21", --0EA8
  X"00", X"40", X"E5", X"C5", X"CD", X"F4", X"0E", X"C1", --0EB0
  X"E1", X"24", X"7C", X"E6", X"07", X"20", X"0A", X"7D", --0EB8
  X"C6", X"20", X"6F", X"3F", X"9F", X"E6", X"F8", X"84", --0EC0
  X"67", X"10", X"E7", X"18", X"0D", X"F3", X"21", X"00", --0EC8
  X"5B", X"06", X"08", X"C5", X"CD", X"F4", X"0E", X"C1", --0ED0
  X"10", X"F9", X"3E", X"04", X"D3", X"FB", X"FB", X"21", --0ED8
  X"00", X"5B", X"FD", X"75", X"46", X"AF", X"47", X"77", --0EE0
  X"23", X"10", X"FC", X"FD", X"CB", X"30", X"8E", X"0E", --0EE8
  X"21", X"C3", X"D9", X"0D", X"78", X"FE", X"03", X"9F", --0EF0
  X"E6", X"02", X"D3", X"FB", X"57", X"CD", X"54", X"1F", --0EF8
  X"38", X"0A", X"3E", X"04", X"D3", X"FB", X"FB", X"CD", --0F00
  X"DF", X"0E", X"CF", X"0C", X"DB", X"FB", X"87", X"F8", --0F08
  X"30", X"EB", X"0E", X"20", X"5E", X"23", X"06", X"08", --0F10
  X"CB", X"12", X"CB", X"13", X"CB", X"1A", X"DB", X"FB", --0F18
  X"1F", X"30", X"FB", X"7A", X"D3", X"FB", X"10", X"F0", --0F20
  X"0D", X"20", X"E9", X"C9", X"2A", X"3D", X"5C", X"E5", --0F28
  X"21", X"7F", X"10", X"E5", X"ED", X"73", X"3D", X"5C", --0F30
  X"CD", X"D4", X"15", X"F5", X"16", X"00", X"FD", X"5E", --0F38
  X"FF", X"21", X"C8", X"00", X"CD", X"B5", X"03", X"F1", --0F40
  X"21", X"38", X"0F", X"E5", X"FE", X"18", X"30", X"31", --0F48
  X"FE", X"07", X"38", X"2D", X"FE", X"10", X"38", X"3A", --0F50
  X"01", X"02", X"00", X"57", X"FE", X"16", X"38", X"0C", --0F58
  X"03", X"FD", X"CB", X"37", X"7E", X"CA", X"1E", X"10", --0F60
  X"CD", X"D4", X"15", X"5F", X"CD", X"D4", X"15", X"D5", --0F68
  X"2A", X"5B", X"5C", X"FD", X"CB", X"07", X"86", X"CD", --0F70
  X"55", X"16", X"C1", X"23", X"70", X"23", X"71", X"18", --0F78
  X"0A", X"FD", X"CB", X"07", X"86", X"2A", X"5B", X"5C", --0F80
  X"CD", X"52", X"16", X"12", X"13", X"ED", X"53", X"5B", --0F88
  X"5C", X"C9", X"5F", X"16", X"00", X"21", X"99", X"0F", --0F90
  X"19", X"5E", X"19", X"E5", X"2A", X"5B", X"5C", X"C9", --0F98
  X"09", X"66", X"6A", X"50", X"B5", X"70", X"7E", X"CF", --0FA0
  X"D4", X"2A", X"49", X"5C", X"FD", X"CB", X"37", X"6E", --0FA8
  X"C2", X"97", X"10", X"CD", X"6E", X"19", X"CD", X"95", --0FB0
  X"16", X"7A", X"B3", X"CA", X"97", X"10", X"E5", X"23", --0FB8
  X"4E", X"23", X"46", X"21", X"0A", X"00", X"09", X"44", --0FC0
  X"4D", X"CD", X"05", X"1F", X"CD", X"97", X"10", X"2A", --0FC8
  X"51", X"5C", X"E3", X"E5", X"3E", X"FF", X"CD", X"01", --0FD0
  X"16", X"E1", X"2B", X"FD", X"35", X"0F", X"CD", X"55", --0FD8
  X"18", X"FD", X"34", X"0F", X"2A", X"59", X"5C", X"23", --0FE0
  X"23", X"23", X"23", X"22", X"5B", X"5C", X"E1", X"CD", --0FE8
  X"15", X"16", X"C9", X"FD", X"CB", X"37", X"6E", X"20", --0FF0
  X"08", X"21", X"49", X"5C", X"CD", X"0F", X"19", X"18", --0FF8
  X"6D", X"FD", X"36", X"00", X"10", X"18", X"1D", X"CD", --1000
  X"31", X"10", X"18", X"05", X"7E", X"FE", X"0D", X"C8", --1008
  X"23", X"22", X"5B", X"5C", X"C9", X"CD", X"31", X"10", --1010
  X"01", X"01", X"00", X"C3", X"E8", X"19", X"CD", X"D4", --1018
  X"15", X"CD", X"D4", X"15", X"E1", X"E1", X"E1", X"22", --1020
  X"3D", X"5C", X"FD", X"CB", X"00", X"7E", X"C0", X"F9", --1028
  X"C9", X"37", X"CD", X"95", X"11", X"ED", X"52", X"19", --1030
  X"23", X"C1", X"D8", X"C5", X"44", X"4D", X"62", X"6B", --1038
  X"23", X"1A", X"E6", X"F0", X"FE", X"10", X"20", X"09", --1040
  X"23", X"1A", X"D6", X"17", X"CE", X"00", X"20", X"01", --1048
  X"23", X"A7", X"ED", X"42", X"09", X"EB", X"38", X"E6", --1050
  X"C9", X"FD", X"CB", X"37", X"6E", X"C0", X"2A", X"49", --1058
  X"5C", X"CD", X"6E", X"19", X"EB", X"CD", X"95", X"16", --1060
  X"21", X"4A", X"5C", X"CD", X"1C", X"19", X"CD", X"95", --1068
  X"17", X"3E", X"00", X"C3", X"01", X"16", X"FD", X"CB", --1070
  X"37", X"7E", X"28", X"A8", X"C3", X"81", X"0F", X"FD", --1078
  X"CB", X"30", X"66", X"28", X"A1", X"FD", X"36", X"00", --1080
  X"FF", X"16", X"00", X"FD", X"5E", X"FE", X"21", X"90", --1088
  X"1A", X"CD", X"B5", X"03", X"C3", X"30", X"0F", X"E5", --1090
  X"CD", X"90", X"11", X"2B", X"CD", X"E5", X"19", X"22", --1098
  X"5B", X"5C", X"FD", X"36", X"07", X"00", X"E1", X"C9", --10A0
  X"FD", X"CB", X"02", X"5E", X"C4", X"1D", X"11", X"A7", --10A8
  X"FD", X"CB", X"01", X"6E", X"C8", X"3A", X"08", X"5C", --10B0
  X"FD", X"CB", X"01", X"AE", X"F5", X"FD", X"CB", X"02", --10B8
  X"6E", X"C4", X"6E", X"0D", X"F1", X"FE", X"20", X"30", --10C0
  X"52", X"FE", X"10", X"30", X"2D", X"FE", X"06", X"30", --10C8
  X"0A", X"47", X"E6", X"01", X"4F", X"78", X"1F", X"C6", --10D0
  X"12", X"18", X"2A", X"20", X"09", X"21", X"6A", X"5C", --10D8
  X"3E", X"08", X"AE", X"77", X"18", X"0E", X"FE", X"0E", --10E0
  X"D8", X"D6", X"0D", X"21", X"41", X"5C", X"BE", X"77", --10E8
  X"20", X"02", X"36", X"00", X"FD", X"CB", X"02", X"DE", --10F0
  X"BF", X"C9", X"47", X"E6", X"07", X"4F", X"3E", X"10", --10F8
  X"CB", X"58", X"20", X"01", X"3C", X"FD", X"71", X"D3", --1100
  X"11", X"0D", X"11", X"18", X"06", X"3A", X"0D", X"5C", --1108
  X"11", X"A8", X"10", X"2A", X"4F", X"5C", X"23", X"23", --1110
  X"73", X"23", X"72", X"37", X"C9", X"CD", X"4D", X"0D", --1118
  X"FD", X"CB", X"02", X"9E", X"FD", X"CB", X"02", X"AE", --1120
  X"2A", X"8A", X"5C", X"E5", X"2A", X"3D", X"5C", X"E5", --1128
  X"21", X"67", X"11", X"E5", X"ED", X"73", X"3D", X"5C", --1130
  X"2A", X"82", X"5C", X"E5", X"37", X"CD", X"95", X"11", --1138
  X"EB", X"CD", X"7D", X"18", X"EB", X"CD", X"E1", X"18", --1140
  X"2A", X"8A", X"5C", X"E3", X"EB", X"CD", X"4D", X"0D", --1148
  X"3A", X"8B", X"5C", X"92", X"38", X"26", X"20", X"06", --1150
  X"7B", X"FD", X"96", X"50", X"30", X"1E", X"3E", X"20", --1158
  X"D5", X"CD", X"F4", X"09", X"D1", X"18", X"E9", X"16", --1160
  X"00", X"FD", X"5E", X"FE", X"21", X"90", X"1A", X"CD", --1168
  X"B5", X"03", X"FD", X"36", X"00", X"FF", X"ED", X"5B", --1170
  X"8A", X"5C", X"18", X"02", X"D1", X"E1", X"E1", X"22", --1178
  X"3D", X"5C", X"C1", X"D5", X"CD", X"D9", X"0D", X"E1", --1180
  X"22", X"82", X"5C", X"FD", X"36", X"26", X"00", X"C9", --1188
  X"2A", X"61", X"5C", X"2B", X"A7", X"ED", X"5B", X"59", --1190
  X"5C", X"FD", X"CB", X"37", X"6E", X"C8", X"ED", X"5B", --1198
  X"61", X"5C", X"D8", X"2A", X"63", X"5C", X"C9", X"7E", --11A0
  X"FE", X"0E", X"01", X"06", X"00", X"CC", X"E8", X"19", --11A8
  X"7E", X"23", X"FE", X"0D", X"20", X"F1", X"C9", X"F3", --11B0
  X"3E", X"FF", X"ED", X"5B", X"B2", X"5C", X"D9", X"ED", --11B8
  X"4B", X"B4", X"5C", X"ED", X"5B", X"38", X"5C", X"2A", --11C0
  X"7B", X"5C", X"D9", X"47", X"3E", X"07", X"D3", X"FE", --11C8
  X"3E", X"3F", X"ED", X"47", X"00", X"00", X"00", X"00", --11D0
  X"00", X"00", X"62", X"6B", X"36", X"02", X"2B", X"BC", --11D8
  X"20", X"FA", X"A7", X"ED", X"52", X"19", X"23", X"30", --11E0
  X"06", X"35", X"28", X"03", X"35", X"28", X"F3", X"2B", --11E8
  X"D9", X"ED", X"43", X"B4", X"5C", X"ED", X"53", X"38", --11F0
  X"5C", X"22", X"7B", X"5C", X"D9", X"04", X"28", X"19", --11F8
  X"22", X"B4", X"5C", X"11", X"AF", X"3E", X"01", X"A8", --1200
  X"00", X"EB", X"ED", X"B8", X"EB", X"23", X"22", X"7B", --1208
  X"5C", X"2B", X"01", X"40", X"00", X"ED", X"43", X"38", --1210
  X"5C", X"22", X"B2", X"5C", X"21", X"00", X"3C", X"22", --1218
  X"36", X"5C", X"2A", X"B2", X"5C", X"36", X"3E", X"2B", --1220
  X"F9", X"2B", X"2B", X"22", X"3D", X"5C", X"ED", X"56", --1228
  X"FD", X"21", X"3A", X"5C", X"FB", X"21", X"B6", X"5C", --1230
  X"22", X"4F", X"5C", X"11", X"AF", X"15", X"01", X"15", --1238
  X"00", X"EB", X"ED", X"B0", X"EB", X"2B", X"22", X"57", --1240
  X"5C", X"23", X"22", X"53", X"5C", X"22", X"4B", X"5C", --1248
  X"36", X"80", X"23", X"22", X"59", X"5C", X"36", X"0D", --1250
  X"23", X"36", X"80", X"23", X"22", X"61", X"5C", X"22", --1258
  X"63", X"5C", X"22", X"65", X"5C", X"3E", X"38", X"32", --1260
  X"8D", X"5C", X"32", X"8F", X"5C", X"32", X"48", X"5C", --1268
  X"21", X"23", X"05", X"22", X"09", X"5C", X"FD", X"35", --1270
  X"C6", X"FD", X"35", X"CA", X"21", X"C6", X"15", X"11", --1278
  X"10", X"5C", X"01", X"0E", X"00", X"ED", X"B0", X"FD", --1280
  X"CB", X"01", X"CE", X"CD", X"DF", X"0E", X"FD", X"36", --1288
  X"31", X"02", X"CD", X"6B", X"0D", X"AF", X"11", X"38", --1290
  X"15", X"CD", X"0A", X"0C", X"FD", X"CB", X"02", X"EE", --1298
  X"18", X"07", X"FD", X"36", X"31", X"02", X"CD", X"95", --12A0
  X"17", X"CD", X"B0", X"16", X"3E", X"00", X"CD", X"01", --12A8
  X"16", X"CD", X"2C", X"0F", X"CD", X"17", X"1B", X"FD", --12B0
  X"CB", X"00", X"7E", X"20", X"12", X"FD", X"CB", X"30", --12B8
  X"66", X"28", X"40", X"2A", X"59", X"5C", X"CD", X"A7", --12C0
  X"11", X"FD", X"36", X"00", X"FF", X"18", X"DD", X"2A", --12C8
  X"59", X"5C", X"22", X"5D", X"5C", X"CD", X"FB", X"19", --12D0
  X"78", X"B1", X"C2", X"5D", X"15", X"DF", X"FE", X"0D", --12D8
  X"28", X"C0", X"FD", X"CB", X"30", X"46", X"C4", X"AF", --12E0
  X"0D", X"CD", X"6E", X"0D", X"3E", X"19", X"FD", X"96", --12E8
  X"4F", X"32", X"8C", X"5C", X"FD", X"CB", X"01", X"FE", --12F0
  X"FD", X"36", X"00", X"FF", X"FD", X"36", X"0A", X"01", --12F8
  X"CD", X"8A", X"1B", X"76", X"FD", X"CB", X"01", X"AE", --1300
  X"FD", X"CB", X"30", X"4E", X"C4", X"CD", X"0E", X"3A", --1308
  X"3A", X"5C", X"3C", X"F5", X"21", X"00", X"00", X"FD", --1310
  X"74", X"37", X"FD", X"74", X"26", X"22", X"0B", X"5C", --1318
  X"21", X"01", X"00", X"22", X"16", X"5C", X"CD", X"B0", --1320
  X"16", X"FD", X"CB", X"37", X"AE", X"CD", X"6E", X"0D", --1328
  X"FD", X"CB", X"02", X"EE", X"F1", X"47", X"FE", X"0A", --1330
  X"38", X"02", X"C6", X"07", X"CD", X"EF", X"15", X"3E", --1338
  X"20", X"D7", X"78", X"11", X"91", X"13", X"CD", X"0A", --1340
  X"0C", X"AF", X"11", X"36", X"15", X"CD", X"0A", X"0C", --1348
  X"ED", X"4B", X"45", X"5C", X"CD", X"1B", X"1A", X"3E", --1350
  X"3A", X"D7", X"FD", X"4E", X"0D", X"06", X"00", X"CD", --1358
  X"1B", X"1A", X"CD", X"97", X"10", X"3A", X"3A", X"5C", --1360
  X"3C", X"28", X"1B", X"FE", X"09", X"28", X"04", X"FE", --1368
  X"15", X"20", X"03", X"FD", X"34", X"0D", X"01", X"03", --1370
  X"00", X"11", X"70", X"5C", X"21", X"44", X"5C", X"CB", --1378
  X"7E", X"28", X"01", X"09", X"ED", X"B8", X"FD", X"36", --1380
  X"0A", X"FF", X"FD", X"CB", X"01", X"9E", X"C3", X"AC", --1388
  X"12", X"80", X"4F", X"CB", X"4E", X"45", X"58", X"54", --1390
  X"20", X"77", X"69", X"74", X"68", X"6F", X"75", X"74", --1398
  X"20", X"46", X"4F", X"D2", X"56", X"61", X"72", X"69", --13A0
  X"61", X"62", X"6C", X"65", X"20", X"6E", X"6F", X"74", --13A8
  X"20", X"66", X"6F", X"75", X"6E", X"E4", X"53", X"75", --13B0
  X"62", X"73", X"63", X"72", X"69", X"70", X"74", X"20", --13B8
  X"77", X"72", X"6F", X"6E", X"E7", X"4F", X"75", X"74", --13C0
  X"20", X"6F", X"66", X"20", X"6D", X"65", X"6D", X"6F", --13C8
  X"72", X"F9", X"4F", X"75", X"74", X"20", X"6F", X"66", --13D0
  X"20", X"73", X"63", X"72", X"65", X"65", X"EE", X"4E", --13D8
  X"75", X"6D", X"62", X"65", X"72", X"20", X"74", X"6F", --13E0
  X"6F", X"20", X"62", X"69", X"E7", X"52", X"45", X"54", --13E8
  X"55", X"52", X"4E", X"20", X"77", X"69", X"74", X"68", --13F0
  X"6F", X"75", X"74", X"20", X"47", X"4F", X"53", X"55", --13F8
  X"C2", X"45", X"6E", X"64", X"20", X"6F", X"66", X"20", --1400
  X"66", X"69", X"6C", X"E5", X"53", X"54", X"4F", X"50", --1408
  X"20", X"73", X"74", X"61", X"74", X"65", X"6D", X"65", --1410
  X"6E", X"F4", X"49", X"6E", X"76", X"61", X"6C", X"69", --1418
  X"64", X"20", X"61", X"72", X"67", X"75", X"6D", X"65", --1420
  X"6E", X"F4", X"49", X"6E", X"74", X"65", X"67", X"65", --1428
  X"72", X"20", X"6F", X"75", X"74", X"20", X"6F", X"66", --1430
  X"20", X"72", X"61", X"6E", X"67", X"E5", X"4E", X"6F", --1438
  X"6E", X"73", X"65", X"6E", X"73", X"65", X"20", X"69", --1440
  X"6E", X"20", X"42", X"41", X"53", X"49", X"C3", X"42", --1448
  X"52", X"45", X"41", X"4B", X"20", X"2D", X"20", X"43", --1450
  X"4F", X"4E", X"54", X"20", X"72", X"65", X"70", X"65", --1458
  X"61", X"74", X"F3", X"4F", X"75", X"74", X"20", X"6F", --1460
  X"66", X"20", X"44", X"41", X"54", X"C1", X"49", X"6E", --1468
  X"76", X"61", X"6C", X"69", X"64", X"20", X"66", X"69", --1470
  X"6C", X"65", X"20", X"6E", X"61", X"6D", X"E5", X"4E", --1478
  X"6F", X"20", X"72", X"6F", X"6F", X"6D", X"20", X"66", --1480
  X"6F", X"72", X"20", X"6C", X"69", X"6E", X"E5", X"53", --1488
  X"54", X"4F", X"50", X"20", X"69", X"6E", X"20", X"49", --1490
  X"4E", X"50", X"55", X"D4", X"46", X"4F", X"52", X"20", --1498
  X"77", X"69", X"74", X"68", X"6F", X"75", X"74", X"20", --14A0
  X"4E", X"45", X"58", X"D4", X"49", X"6E", X"76", X"61", --14A8
  X"6C", X"69", X"64", X"20", X"49", X"2F", X"4F", X"20", --14B0
  X"64", X"65", X"76", X"69", X"63", X"E5", X"49", X"6E", --14B8
  X"76", X"61", X"6C", X"69", X"64", X"20", X"63", X"6F", --14C0
  X"6C", X"6F", X"75", X"F2", X"42", X"52", X"45", X"41", --14C8
  X"4B", X"20", X"69", X"6E", X"74", X"6F", X"20", X"70", --14D0
  X"72", X"6F", X"67", X"72", X"61", X"ED", X"52", X"41", --14D8
  X"4D", X"54", X"4F", X"50", X"20", X"6E", X"6F", X"20", --14E0
  X"67", X"6F", X"6F", X"E4", X"53", X"74", X"61", X"74", --14E8
  X"65", X"6D", X"65", X"6E", X"74", X"20", X"6C", X"6F", --14F0
  X"73", X"F4", X"49", X"6E", X"76", X"61", X"6C", X"69", --14F8
  X"64", X"20", X"73", X"74", X"72", X"65", X"61", X"ED", --1500
  X"46", X"4E", X"20", X"77", X"69", X"74", X"68", X"6F", --1508
  X"75", X"74", X"20", X"44", X"45", X"C6", X"50", X"61", --1510
  X"72", X"61", X"6D", X"65", X"74", X"65", X"72", X"20", --1518
  X"65", X"72", X"72", X"6F", X"F2", X"54", X"61", X"70", --1520
  X"65", X"20", X"6C", X"6F", X"61", X"64", X"69", X"6E", --1528
  X"67", X"20", X"65", X"72", X"72", X"6F", X"F2", X"2C", --1530
  X"A0", X"7F", X"20", X"31", X"39", X"38", X"32", X"20", --1538
  X"53", X"69", X"6E", X"63", X"6C", X"61", X"69", X"72", --1540
  X"20", X"52", X"65", X"73", X"65", X"61", X"72", X"63", --1548
  X"68", X"20", X"4C", X"74", X"E4", X"3E", X"10", X"01", --1550
  X"00", X"00", X"C3", X"13", X"13", X"ED", X"43", X"49", --1558
  X"5C", X"2A", X"5D", X"5C", X"EB", X"21", X"55", X"15", --1560
  X"E5", X"2A", X"61", X"5C", X"37", X"ED", X"52", X"E5", --1568
  X"60", X"69", X"CD", X"6E", X"19", X"20", X"06", X"CD", --1570
  X"B8", X"19", X"CD", X"E8", X"19", X"C1", X"79", X"3D", --1578
  X"B0", X"28", X"28", X"C5", X"03", X"03", X"03", X"03", --1580
  X"2B", X"ED", X"5B", X"53", X"5C", X"D5", X"CD", X"55", --1588
  X"16", X"E1", X"22", X"53", X"5C", X"C1", X"C5", X"13", --1590
  X"2A", X"61", X"5C", X"2B", X"2B", X"ED", X"B8", X"2A", --1598
  X"49", X"5C", X"EB", X"C1", X"70", X"2B", X"71", X"2B", --15A0
  X"73", X"2B", X"72", X"F1", X"C3", X"A2", X"12", X"F4", --15A8
  X"09", X"A8", X"10", X"4B", X"F4", X"09", X"C4", X"15", --15B0
  X"53", X"81", X"0F", X"C4", X"15", X"52", X"F4", X"09", --15B8
  X"C4", X"15", X"50", X"80", X"CF", X"12", X"01", X"00", --15C0
  X"06", X"00", X"0B", X"00", X"01", X"00", X"01", X"00", --15C8
  X"06", X"00", X"10", X"00", X"FD", X"CB", X"02", X"6E", --15D0
  X"20", X"04", X"FD", X"CB", X"02", X"DE", X"CD", X"E6", --15D8
  X"15", X"D8", X"28", X"FA", X"CF", X"07", X"D9", X"E5", --15E0
  X"2A", X"51", X"5C", X"23", X"23", X"18", X"08", X"1E", --15E8
  X"30", X"83", X"D9", X"E5", X"2A", X"51", X"5C", X"5E", --15F0
  X"23", X"56", X"EB", X"CD", X"2C", X"16", X"E1", X"D9", --15F8
  X"C9", X"87", X"C6", X"16", X"6F", X"26", X"5C", X"5E", --1600
  X"23", X"56", X"7A", X"B3", X"20", X"02", X"CF", X"17", --1608
  X"1B", X"2A", X"4F", X"5C", X"19", X"22", X"51", X"5C", --1610
  X"FD", X"CB", X"30", X"A6", X"23", X"23", X"23", X"23", --1618
  X"4E", X"21", X"2D", X"16", X"CD", X"DC", X"16", X"D0", --1620
  X"16", X"00", X"5E", X"19", X"E9", X"4B", X"06", X"53", --1628
  X"12", X"50", X"1B", X"00", X"FD", X"CB", X"02", X"C6", --1630
  X"FD", X"CB", X"01", X"AE", X"FD", X"CB", X"30", X"E6", --1638
  X"18", X"04", X"FD", X"CB", X"02", X"86", X"FD", X"CB", --1640
  X"01", X"8E", X"C3", X"4D", X"0D", X"FD", X"CB", X"01", --1648
  X"CE", X"C9", X"01", X"01", X"00", X"E5", X"CD", X"05", --1650
  X"1F", X"E1", X"CD", X"64", X"16", X"2A", X"65", X"5C", --1658
  X"EB", X"ED", X"B8", X"C9", X"F5", X"E5", X"21", X"4B", --1660
  X"5C", X"3E", X"0E", X"5E", X"23", X"56", X"E3", X"A7", --1668
  X"ED", X"52", X"19", X"E3", X"30", X"09", X"D5", X"EB", --1670
  X"09", X"EB", X"72", X"2B", X"73", X"23", X"D1", X"23", --1678
  X"3D", X"20", X"E8", X"EB", X"D1", X"F1", X"A7", X"ED", --1680
  X"52", X"44", X"4D", X"03", X"19", X"EB", X"C9", X"00", --1688
  X"00", X"EB", X"11", X"8F", X"16", X"7E", X"E6", X"C0", --1690
  X"20", X"F7", X"56", X"23", X"5E", X"C9", X"2A", X"63", --1698
  X"5C", X"2B", X"CD", X"55", X"16", X"23", X"23", X"C1", --16A0
  X"ED", X"43", X"61", X"5C", X"C1", X"EB", X"23", X"C9", --16A8
  X"2A", X"59", X"5C", X"36", X"0D", X"22", X"5B", X"5C", --16B0
  X"23", X"36", X"80", X"23", X"22", X"61", X"5C", X"2A", --16B8
  X"61", X"5C", X"22", X"63", X"5C", X"2A", X"63", X"5C", --16C0
  X"22", X"65", X"5C", X"E5", X"21", X"92", X"5C", X"22", --16C8
  X"68", X"5C", X"E1", X"C9", X"ED", X"5B", X"59", X"5C", --16D0
  X"C3", X"E5", X"19", X"23", X"7E", X"A7", X"C8", X"B9", --16D8
  X"23", X"20", X"F8", X"37", X"C9", X"CD", X"1E", X"17", --16E0
  X"CD", X"01", X"17", X"01", X"00", X"00", X"11", X"E2", --16E8
  X"A3", X"EB", X"19", X"38", X"07", X"01", X"D4", X"15", --16F0
  X"09", X"4E", X"23", X"46", X"EB", X"71", X"23", X"70", --16F8
  X"C9", X"E5", X"2A", X"4F", X"5C", X"09", X"23", X"23", --1700
  X"23", X"4E", X"EB", X"21", X"16", X"17", X"CD", X"DC", --1708
  X"16", X"4E", X"06", X"00", X"09", X"E9", X"4B", X"05", --1710
  X"53", X"03", X"50", X"01", X"E1", X"C9", X"CD", X"94", --1718
  X"1E", X"FE", X"10", X"38", X"02", X"CF", X"17", X"C6", --1720
  X"03", X"07", X"21", X"10", X"5C", X"4F", X"06", X"00", --1728
  X"09", X"4E", X"23", X"46", X"2B", X"C9", X"EF", X"01", --1730
  X"38", X"CD", X"1E", X"17", X"78", X"B1", X"28", X"16", --1738
  X"EB", X"2A", X"4F", X"5C", X"09", X"23", X"23", X"23", --1740
  X"7E", X"EB", X"FE", X"4B", X"28", X"08", X"FE", X"53", --1748
  X"28", X"04", X"FE", X"50", X"20", X"CF", X"CD", X"5D", --1750
  X"17", X"73", X"23", X"72", X"C9", X"E5", X"CD", X"F1", --1758
  X"2B", X"78", X"B1", X"20", X"02", X"CF", X"0E", X"C5", --1760
  X"1A", X"E6", X"DF", X"4F", X"21", X"7A", X"17", X"CD", --1768
  X"DC", X"16", X"30", X"F1", X"4E", X"06", X"00", X"09", --1770
  X"C1", X"E9", X"4B", X"06", X"53", X"08", X"50", X"0A", --1778
  X"00", X"1E", X"01", X"18", X"06", X"1E", X"06", X"18", --1780
  X"02", X"1E", X"10", X"0B", X"78", X"B1", X"20", X"D5", --1788
  X"57", X"E1", X"C9", X"18", X"90", X"ED", X"73", X"3F", --1790
  X"5C", X"FD", X"36", X"02", X"10", X"CD", X"AF", X"0D", --1798
  X"FD", X"CB", X"02", X"C6", X"FD", X"46", X"31", X"CD", --17A0
  X"44", X"0E", X"FD", X"CB", X"02", X"86", X"FD", X"CB", --17A8
  X"30", X"C6", X"2A", X"49", X"5C", X"ED", X"5B", X"6C", --17B0
  X"5C", X"A7", X"ED", X"52", X"19", X"38", X"22", X"D5", --17B8
  X"CD", X"6E", X"19", X"11", X"C0", X"02", X"EB", X"ED", --17C0
  X"52", X"E3", X"CD", X"6E", X"19", X"C1", X"C5", X"CD", --17C8
  X"B8", X"19", X"C1", X"09", X"38", X"0E", X"EB", X"56", --17D0
  X"23", X"5E", X"2B", X"ED", X"53", X"6C", X"5C", X"18", --17D8
  X"ED", X"22", X"6C", X"5C", X"2A", X"6C", X"5C", X"CD", --17E0
  X"6E", X"19", X"28", X"01", X"EB", X"CD", X"33", X"18", --17E8
  X"FD", X"CB", X"02", X"A6", X"C9", X"3E", X"03", X"18", --17F0
  X"02", X"3E", X"02", X"FD", X"36", X"02", X"00", X"CD", --17F8
  X"30", X"25", X"C4", X"01", X"16", X"DF", X"CD", X"70", --1800
  X"20", X"38", X"14", X"DF", X"FE", X"3B", X"28", X"04", --1808
  X"FE", X"2C", X"20", X"06", X"E7", X"CD", X"82", X"1C", --1810
  X"18", X"08", X"CD", X"E6", X"1C", X"18", X"03", X"CD", --1818
  X"DE", X"1C", X"CD", X"EE", X"1B", X"CD", X"99", X"1E", --1820
  X"78", X"E6", X"3F", X"67", X"69", X"22", X"49", X"5C", --1828
  X"CD", X"6E", X"19", X"1E", X"01", X"CD", X"55", X"18", --1830
  X"D7", X"FD", X"CB", X"02", X"66", X"28", X"F6", X"3A", --1838
  X"6B", X"5C", X"FD", X"96", X"4F", X"20", X"EE", X"AB", --1840
  X"C8", X"E5", X"D5", X"21", X"6C", X"5C", X"CD", X"0F", --1848
  X"19", X"D1", X"E1", X"18", X"E0", X"ED", X"4B", X"49", --1850
  X"5C", X"CD", X"80", X"19", X"16", X"3E", X"28", X"05", --1858
  X"11", X"00", X"00", X"CB", X"13", X"FD", X"73", X"2D", --1860
  X"7E", X"FE", X"40", X"C1", X"D0", X"C5", X"CD", X"28", --1868
  X"1A", X"23", X"23", X"23", X"FD", X"CB", X"01", X"86", --1870
  X"7A", X"A7", X"28", X"05", X"D7", X"FD", X"CB", X"01", --1878
  X"C6", X"D5", X"EB", X"FD", X"CB", X"30", X"96", X"21", --1880
  X"3B", X"5C", X"CB", X"96", X"FD", X"CB", X"37", X"6E", --1888
  X"28", X"02", X"CB", X"D6", X"2A", X"5F", X"5C", X"A7", --1890
  X"ED", X"52", X"20", X"05", X"3E", X"3F", X"CD", X"C1", --1898
  X"18", X"CD", X"E1", X"18", X"EB", X"7E", X"CD", X"B6", --18A0
  X"18", X"23", X"FE", X"0D", X"28", X"06", X"EB", X"CD", --18A8
  X"37", X"19", X"18", X"E0", X"D1", X"C9", X"FE", X"0E", --18B0
  X"C0", X"23", X"23", X"23", X"23", X"23", X"23", X"7E", --18B8
  X"C9", X"D9", X"2A", X"8F", X"5C", X"E5", X"CB", X"BC", --18C0
  X"CB", X"FD", X"22", X"8F", X"5C", X"21", X"91", X"5C", --18C8
  X"56", X"D5", X"36", X"00", X"CD", X"F4", X"09", X"E1", --18D0
  X"FD", X"74", X"57", X"E1", X"22", X"8F", X"5C", X"D9", --18D8
  X"C9", X"2A", X"5B", X"5C", X"A7", X"ED", X"52", X"C0", --18E0
  X"3A", X"41", X"5C", X"CB", X"07", X"28", X"04", X"C6", --18E8
  X"43", X"18", X"16", X"21", X"3B", X"5C", X"CB", X"9E", --18F0
  X"3E", X"4B", X"CB", X"56", X"28", X"0B", X"CB", X"DE", --18F8
  X"3C", X"FD", X"CB", X"30", X"5E", X"28", X"02", X"3E", --1900
  X"43", X"D5", X"CD", X"C1", X"18", X"D1", X"C9", X"5E", --1908
  X"23", X"56", X"E5", X"EB", X"23", X"CD", X"6E", X"19", --1910
  X"CD", X"95", X"16", X"E1", X"FD", X"CB", X"37", X"6E", --1918
  X"C0", X"72", X"2B", X"73", X"C9", X"7B", X"A7", X"F8", --1920
  X"18", X"0D", X"AF", X"09", X"3C", X"38", X"FC", X"ED", --1928
  X"42", X"3D", X"28", X"F1", X"C3", X"EF", X"15", X"CD", --1930
  X"1B", X"2D", X"30", X"30", X"FE", X"21", X"38", X"2C", --1938
  X"FD", X"CB", X"01", X"96", X"FE", X"CB", X"28", X"24", --1940
  X"FE", X"3A", X"20", X"0E", X"FD", X"CB", X"37", X"6E", --1948
  X"20", X"16", X"FD", X"CB", X"30", X"56", X"28", X"14", --1950
  X"18", X"0E", X"FE", X"22", X"20", X"0A", X"F5", X"3A", --1958
  X"6A", X"5C", X"EE", X"04", X"32", X"6A", X"5C", X"F1", --1960
  X"FD", X"CB", X"01", X"D6", X"D7", X"C9", X"E5", X"2A", --1968
  X"53", X"5C", X"54", X"5D", X"C1", X"CD", X"80", X"19", --1970
  X"D0", X"C5", X"CD", X"B8", X"19", X"EB", X"18", X"F4", --1978
  X"7E", X"B8", X"C0", X"23", X"7E", X"2B", X"B9", X"C9", --1980
  X"23", X"23", X"23", X"22", X"5D", X"5C", X"0E", X"00", --1988
  X"15", X"C8", X"E7", X"BB", X"20", X"04", X"A7", X"C9", --1990
  X"23", X"7E", X"CD", X"B6", X"18", X"22", X"5D", X"5C", --1998
  X"FE", X"22", X"20", X"01", X"0D", X"FE", X"3A", X"28", --19A0
  X"04", X"FE", X"CB", X"20", X"04", X"CB", X"41", X"28", --19A8
  X"DF", X"FE", X"0D", X"20", X"E3", X"15", X"37", X"C9", --19B0
  X"E5", X"7E", X"FE", X"40", X"38", X"17", X"CB", X"6F", --19B8
  X"28", X"14", X"87", X"FA", X"C7", X"19", X"3F", X"01", --19C0
  X"05", X"00", X"30", X"02", X"0E", X"12", X"17", X"23", --19C8
  X"7E", X"30", X"FB", X"18", X"06", X"23", X"23", X"4E", --19D0
  X"23", X"46", X"23", X"09", X"D1", X"A7", X"ED", X"52", --19D8
  X"44", X"4D", X"19", X"EB", X"C9", X"CD", X"DD", X"19", --19E0
  X"C5", X"78", X"2F", X"47", X"79", X"2F", X"4F", X"03", --19E8
  X"CD", X"64", X"16", X"EB", X"E1", X"19", X"D5", X"ED", --19F0
  X"B0", X"E1", X"C9", X"2A", X"59", X"5C", X"2B", X"22", --19F8
  X"5D", X"5C", X"E7", X"21", X"92", X"5C", X"22", X"65", --1A00
  X"5C", X"CD", X"3B", X"2D", X"CD", X"A2", X"2D", X"38", --1A08
  X"04", X"21", X"F0", X"D8", X"09", X"DA", X"8A", X"1C", --1A10
  X"C3", X"C5", X"16", X"D5", X"E5", X"AF", X"CB", X"78", --1A18
  X"20", X"20", X"60", X"69", X"1E", X"FF", X"18", X"08", --1A20
  X"D5", X"56", X"23", X"5E", X"E5", X"EB", X"1E", X"20", --1A28
  X"01", X"18", X"FC", X"CD", X"2A", X"19", X"01", X"9C", --1A30
  X"FF", X"CD", X"2A", X"19", X"0E", X"F6", X"CD", X"2A", --1A38
  X"19", X"7D", X"CD", X"EF", X"15", X"E1", X"D1", X"C9", --1A40
  X"B1", X"CB", X"BC", X"BF", X"C4", X"AF", X"B4", X"93", --1A48
  X"91", X"92", X"95", X"98", X"98", X"98", X"98", X"98", --1A50
  X"98", X"98", X"7F", X"81", X"2E", X"6C", X"6E", X"70", --1A58
  X"48", X"94", X"56", X"3F", X"41", X"2B", X"17", X"1F", --1A60
  X"37", X"77", X"44", X"0F", X"59", X"2B", X"43", X"2D", --1A68
  X"51", X"3A", X"6D", X"42", X"0D", X"49", X"5C", X"44", --1A70
  X"15", X"5D", X"01", X"3D", X"02", X"06", X"00", X"67", --1A78
  X"1E", X"06", X"CB", X"05", X"F0", X"1C", X"06", X"00", --1A80
  X"ED", X"1E", X"00", X"EE", X"1C", X"00", X"23", X"1F", --1A88
  X"04", X"3D", X"06", X"CC", X"06", X"05", X"03", X"1D", --1A90
  X"04", X"00", X"AB", X"1D", X"05", X"CD", X"1F", X"05", --1A98
  X"89", X"20", X"05", X"02", X"2C", X"05", X"B2", X"1B", --1AA0
  X"00", X"B7", X"11", X"03", X"A1", X"1E", X"05", X"F9", --1AA8
  X"17", X"08", X"00", X"80", X"1E", X"03", X"4F", X"1E", --1AB0
  X"00", X"5F", X"1E", X"03", X"AC", X"1E", X"00", X"6B", --1AB8
  X"0D", X"09", X"00", X"DC", X"22", X"06", X"00", X"3A", --1AC0
  X"1F", X"05", X"ED", X"1D", X"05", X"27", X"1E", X"03", --1AC8
  X"42", X"1E", X"09", X"05", X"82", X"23", X"00", X"AC", --1AD0
  X"0E", X"05", X"C9", X"1F", X"05", X"F5", X"17", X"0B", --1AD8
  X"0B", X"0B", X"0B", X"08", X"00", X"F8", X"03", X"09", --1AE0
  X"05", X"20", X"23", X"07", X"07", X"07", X"07", X"07", --1AE8
  X"07", X"08", X"00", X"7A", X"1E", X"06", X"00", X"94", --1AF0
  X"22", X"05", X"60", X"1F", X"06", X"2C", X"0A", X"00", --1AF8
  X"36", X"17", X"06", X"00", X"E5", X"16", X"0A", X"00", --1B00
  X"93", X"17", X"0A", X"2C", X"0A", X"00", X"93", X"17", --1B08
  X"0A", X"00", X"93", X"17", X"00", X"93", X"17", X"FD", --1B10
  X"CB", X"01", X"BE", X"CD", X"FB", X"19", X"AF", X"32", --1B18
  X"47", X"5C", X"3D", X"32", X"3A", X"5C", X"18", X"01", --1B20
  X"E7", X"CD", X"BF", X"16", X"FD", X"34", X"0D", X"FA", --1B28
  X"8A", X"1C", X"DF", X"06", X"00", X"FE", X"0D", X"28", --1B30
  X"7A", X"FE", X"3A", X"28", X"EB", X"21", X"76", X"1B", --1B38
  X"E5", X"4F", X"E7", X"79", X"D6", X"CE", X"DA", X"8A", --1B40
  X"1C", X"4F", X"21", X"48", X"1A", X"09", X"4E", X"09", --1B48
  X"18", X"03", X"2A", X"74", X"5C", X"7E", X"23", X"22", --1B50
  X"74", X"5C", X"01", X"52", X"1B", X"C5", X"4F", X"FE", --1B58
  X"20", X"30", X"0C", X"21", X"01", X"1C", X"06", X"00", --1B60
  X"09", X"4E", X"09", X"E5", X"DF", X"05", X"C9", X"DF", --1B68
  X"B9", X"C2", X"8A", X"1C", X"E7", X"C9", X"CD", X"54", --1B70
  X"1F", X"38", X"02", X"CF", X"14", X"FD", X"CB", X"0A", --1B78
  X"7E", X"20", X"71", X"2A", X"42", X"5C", X"CB", X"7C", --1B80
  X"28", X"14", X"21", X"FE", X"FF", X"22", X"45", X"5C", --1B88
  X"2A", X"61", X"5C", X"2B", X"ED", X"5B", X"59", X"5C", --1B90
  X"1B", X"3A", X"44", X"5C", X"18", X"33", X"CD", X"6E", --1B98
  X"19", X"3A", X"44", X"5C", X"28", X"19", X"A7", X"20", --1BA0
  X"43", X"47", X"7E", X"E6", X"C0", X"78", X"28", X"0F", --1BA8
  X"CF", X"FF", X"C1", X"CD", X"30", X"25", X"C8", X"2A", --1BB0
  X"55", X"5C", X"3E", X"C0", X"A6", X"C0", X"AF", X"FE", --1BB8
  X"01", X"CE", X"00", X"56", X"23", X"5E", X"ED", X"53", --1BC0
  X"45", X"5C", X"23", X"5E", X"23", X"56", X"EB", X"19", --1BC8
  X"23", X"22", X"55", X"5C", X"EB", X"22", X"5D", X"5C", --1BD0
  X"57", X"1E", X"00", X"FD", X"36", X"0A", X"FF", X"15", --1BD8
  X"FD", X"72", X"0D", X"CA", X"28", X"1B", X"14", X"CD", --1BE0
  X"8B", X"19", X"28", X"08", X"CF", X"16", X"CD", X"30", --1BE8
  X"25", X"C0", X"C1", X"C1", X"DF", X"FE", X"0D", X"28", --1BF0
  X"BA", X"FE", X"3A", X"CA", X"28", X"1B", X"C3", X"8A", --1BF8
  X"1C", X"0F", X"1D", X"4B", X"09", X"67", X"0B", X"7B", --1C00
  X"8E", X"71", X"B4", X"81", X"CF", X"CD", X"DE", X"1C", --1C08
  X"BF", X"C1", X"CC", X"EE", X"1B", X"EB", X"2A", X"74", --1C10
  X"5C", X"4E", X"23", X"46", X"EB", X"C5", X"C9", X"CD", --1C18
  X"B2", X"28", X"FD", X"36", X"37", X"00", X"30", X"08", --1C20
  X"FD", X"CB", X"37", X"CE", X"20", X"18", X"CF", X"01", --1C28
  X"CC", X"96", X"29", X"FD", X"CB", X"01", X"76", X"20", --1C30
  X"0D", X"AF", X"CD", X"30", X"25", X"C4", X"F1", X"2B", --1C38
  X"21", X"71", X"5C", X"B6", X"77", X"EB", X"ED", X"43", --1C40
  X"72", X"5C", X"22", X"4D", X"5C", X"C9", X"C1", X"CD", --1C48
  X"56", X"1C", X"CD", X"EE", X"1B", X"C9", X"3A", X"3B", --1C50
  X"5C", X"F5", X"CD", X"FB", X"24", X"F1", X"FD", X"56", --1C58
  X"01", X"AA", X"E6", X"40", X"20", X"24", X"CB", X"7A", --1C60
  X"C2", X"FF", X"2A", X"C9", X"CD", X"B2", X"28", X"F5", --1C68
  X"79", X"F6", X"9F", X"3C", X"20", X"14", X"F1", X"18", --1C70
  X"A9", X"E7", X"CD", X"82", X"1C", X"FE", X"2C", X"20", --1C78
  X"09", X"E7", X"CD", X"FB", X"24", X"FD", X"CB", X"01", --1C80
  X"76", X"C0", X"CF", X"0B", X"CD", X"FB", X"24", X"FD", --1C88
  X"CB", X"01", X"76", X"C8", X"18", X"F4", X"FD", X"CB", --1C90
  X"01", X"7E", X"FD", X"CB", X"02", X"86", X"C4", X"4D", --1C98
  X"0D", X"F1", X"3A", X"74", X"5C", X"D6", X"13", X"CD", --1CA0
  X"FC", X"21", X"CD", X"EE", X"1B", X"2A", X"8F", X"5C", --1CA8
  X"22", X"8D", X"5C", X"21", X"91", X"5C", X"7E", X"07", --1CB0
  X"AE", X"E6", X"AA", X"AE", X"77", X"C9", X"CD", X"30", --1CB8
  X"25", X"28", X"13", X"FD", X"CB", X"02", X"86", X"CD", --1CC0
  X"4D", X"0D", X"21", X"90", X"5C", X"7E", X"F6", X"F8", --1CC8
  X"77", X"FD", X"CB", X"57", X"B6", X"DF", X"CD", X"E2", --1CD0
  X"21", X"18", X"9F", X"C3", X"05", X"06", X"FE", X"0D", --1CD8
  X"28", X"04", X"FE", X"3A", X"20", X"9C", X"CD", X"30", --1CE0
  X"25", X"C8", X"EF", X"A0", X"38", X"C9", X"CF", X"08", --1CE8
  X"C1", X"CD", X"30", X"25", X"28", X"0A", X"EF", X"02", --1CF0
  X"38", X"EB", X"CD", X"E9", X"34", X"DA", X"B3", X"1B", --1CF8
  X"C3", X"29", X"1B", X"FE", X"CD", X"20", X"09", X"E7", --1D00
  X"CD", X"82", X"1C", X"CD", X"EE", X"1B", X"18", X"06", --1D08
  X"CD", X"EE", X"1B", X"EF", X"A1", X"38", X"EF", X"C0", --1D10
  X"02", X"01", X"E0", X"01", X"38", X"CD", X"FF", X"2A", --1D18
  X"22", X"68", X"5C", X"2B", X"7E", X"CB", X"FE", X"01", --1D20
  X"06", X"00", X"09", X"07", X"38", X"06", X"0E", X"0D", --1D28
  X"CD", X"55", X"16", X"23", X"E5", X"EF", X"02", X"02", --1D30
  X"38", X"E1", X"EB", X"0E", X"0A", X"ED", X"B0", X"2A", --1D38
  X"45", X"5C", X"EB", X"73", X"23", X"72", X"FD", X"56", --1D40
  X"0D", X"14", X"23", X"72", X"CD", X"DA", X"1D", X"D0", --1D48
  X"FD", X"46", X"38", X"2A", X"45", X"5C", X"22", X"42", --1D50
  X"5C", X"3A", X"47", X"5C", X"ED", X"44", X"57", X"2A", --1D58
  X"5D", X"5C", X"1E", X"F3", X"C5", X"ED", X"4B", X"55", --1D60
  X"5C", X"CD", X"86", X"1D", X"ED", X"43", X"55", X"5C", --1D68
  X"C1", X"38", X"11", X"E7", X"F6", X"20", X"B8", X"28", --1D70
  X"03", X"E7", X"18", X"E8", X"E7", X"3E", X"01", X"92", --1D78
  X"32", X"44", X"5C", X"C9", X"CF", X"11", X"7E", X"FE", --1D80
  X"3A", X"28", X"18", X"23", X"7E", X"E6", X"C0", X"37", --1D88
  X"C0", X"46", X"23", X"4E", X"ED", X"43", X"42", X"5C", --1D90
  X"23", X"4E", X"23", X"46", X"E5", X"09", X"44", X"4D", --1D98
  X"E1", X"16", X"00", X"C5", X"CD", X"8B", X"19", X"C1", --1DA0
  X"D0", X"18", X"E0", X"FD", X"CB", X"37", X"4E", X"C2", --1DA8
  X"2E", X"1C", X"2A", X"4D", X"5C", X"CB", X"7E", X"28", --1DB0
  X"1F", X"23", X"22", X"68", X"5C", X"EF", X"E0", X"E2", --1DB8
  X"0F", X"C0", X"02", X"38", X"CD", X"DA", X"1D", X"D8", --1DC0
  X"2A", X"68", X"5C", X"11", X"0F", X"00", X"19", X"5E", --1DC8
  X"23", X"56", X"23", X"66", X"EB", X"C3", X"73", X"1E", --1DD0
  X"CF", X"00", X"EF", X"E1", X"E0", X"E2", X"36", X"00", --1DD8
  X"02", X"01", X"03", X"37", X"00", X"04", X"38", X"A7", --1DE0
  X"C9", X"38", X"37", X"C9", X"E7", X"CD", X"1F", X"1C", --1DE8
  X"CD", X"30", X"25", X"28", X"29", X"DF", X"22", X"5F", --1DF0
  X"5C", X"2A", X"57", X"5C", X"7E", X"FE", X"2C", X"28", --1DF8
  X"09", X"1E", X"E4", X"CD", X"86", X"1D", X"30", X"02", --1E00
  X"CF", X"0D", X"CD", X"77", X"00", X"CD", X"56", X"1C", --1E08
  X"DF", X"22", X"57", X"5C", X"2A", X"5F", X"5C", X"FD", --1E10
  X"36", X"26", X"00", X"CD", X"78", X"00", X"DF", X"FE", --1E18
  X"2C", X"28", X"C9", X"CD", X"EE", X"1B", X"C9", X"CD", --1E20
  X"30", X"25", X"20", X"0B", X"CD", X"FB", X"24", X"FE", --1E28
  X"2C", X"C4", X"EE", X"1B", X"E7", X"18", X"F5", X"3E", --1E30
  X"E4", X"47", X"ED", X"B9", X"11", X"00", X"02", X"C3", --1E38
  X"8B", X"19", X"CD", X"99", X"1E", X"60", X"69", X"CD", --1E40
  X"6E", X"19", X"2B", X"22", X"57", X"5C", X"C9", X"CD", --1E48
  X"99", X"1E", X"78", X"B1", X"20", X"04", X"ED", X"4B", --1E50
  X"78", X"5C", X"ED", X"43", X"76", X"5C", X"C9", X"2A", --1E58
  X"6E", X"5C", X"FD", X"56", X"36", X"18", X"0C", X"CD", --1E60
  X"99", X"1E", X"60", X"69", X"16", X"00", X"7C", X"FE", --1E68
  X"F0", X"30", X"2C", X"22", X"42", X"5C", X"FD", X"72", --1E70
  X"0A", X"C9", X"CD", X"85", X"1E", X"ED", X"79", X"C9", --1E78
  X"CD", X"85", X"1E", X"02", X"C9", X"CD", X"D5", X"2D", --1E80
  X"38", X"15", X"28", X"02", X"ED", X"44", X"F5", X"CD", --1E88
  X"99", X"1E", X"F1", X"C9", X"CD", X"D5", X"2D", X"18", --1E90
  X"03", X"CD", X"A2", X"2D", X"38", X"01", X"C8", X"CF", --1E98
  X"0A", X"CD", X"67", X"1E", X"01", X"00", X"00", X"CD", --1EA0
  X"45", X"1E", X"18", X"03", X"CD", X"99", X"1E", X"78", --1EA8
  X"B1", X"20", X"04", X"ED", X"4B", X"B2", X"5C", X"C5", --1EB0
  X"ED", X"5B", X"4B", X"5C", X"2A", X"59", X"5C", X"2B", --1EB8
  X"CD", X"E5", X"19", X"CD", X"6B", X"0D", X"2A", X"65", --1EC0
  X"5C", X"11", X"32", X"00", X"19", X"D1", X"ED", X"52", --1EC8
  X"30", X"08", X"2A", X"B4", X"5C", X"A7", X"ED", X"52", --1ED0
  X"30", X"02", X"CF", X"15", X"EB", X"22", X"B2", X"5C", --1ED8
  X"D1", X"C1", X"36", X"3E", X"2B", X"F9", X"C5", X"ED", --1EE0
  X"73", X"3D", X"5C", X"EB", X"E9", X"D1", X"FD", X"66", --1EE8
  X"0D", X"24", X"E3", X"33", X"ED", X"4B", X"45", X"5C", --1EF0
  X"C5", X"E5", X"ED", X"73", X"3D", X"5C", X"D5", X"CD", --1EF8
  X"67", X"1E", X"01", X"14", X"00", X"2A", X"65", X"5C", --1F00
  X"09", X"38", X"0A", X"EB", X"21", X"50", X"00", X"19", --1F08
  X"38", X"03", X"ED", X"72", X"D8", X"2E", X"03", X"C3", --1F10
  X"55", X"00", X"01", X"00", X"00", X"CD", X"05", X"1F", --1F18
  X"44", X"4D", X"C9", X"C1", X"E1", X"D1", X"7A", X"FE", --1F20
  X"3E", X"28", X"0B", X"3B", X"E3", X"EB", X"ED", X"73", --1F28
  X"3D", X"5C", X"C5", X"C3", X"73", X"1E", X"D5", X"E5", --1F30
  X"CF", X"06", X"CD", X"99", X"1E", X"76", X"0B", X"78", --1F38
  X"B1", X"28", X"0C", X"78", X"A1", X"3C", X"20", X"01", --1F40
  X"03", X"FD", X"CB", X"01", X"6E", X"28", X"EE", X"FD", --1F48
  X"CB", X"01", X"AE", X"C9", X"3E", X"7F", X"DB", X"FE", --1F50
  X"1F", X"D8", X"3E", X"FE", X"DB", X"FE", X"1F", X"C9", --1F58
  X"CD", X"30", X"25", X"28", X"05", X"3E", X"CE", X"C3", --1F60
  X"39", X"1E", X"FD", X"CB", X"01", X"F6", X"CD", X"8D", --1F68
  X"2C", X"30", X"16", X"E7", X"FE", X"24", X"20", X"05", --1F70
  X"FD", X"CB", X"01", X"B6", X"E7", X"FE", X"28", X"20", --1F78
  X"3C", X"E7", X"FE", X"29", X"28", X"20", X"CD", X"8D", --1F80
  X"2C", X"D2", X"8A", X"1C", X"EB", X"E7", X"FE", X"24", --1F88
  X"20", X"02", X"EB", X"E7", X"EB", X"01", X"06", X"00", --1F90
  X"CD", X"55", X"16", X"23", X"23", X"36", X"0E", X"FE", --1F98
  X"2C", X"20", X"03", X"E7", X"18", X"E0", X"FE", X"29", --1FA0
  X"20", X"13", X"E7", X"FE", X"3D", X"20", X"0E", X"E7", --1FA8
  X"3A", X"3B", X"5C", X"F5", X"CD", X"FB", X"24", X"F1", --1FB0
  X"FD", X"AE", X"01", X"E6", X"40", X"C2", X"8A", X"1C", --1FB8
  X"CD", X"EE", X"1B", X"CD", X"30", X"25", X"E1", X"C8", --1FC0
  X"E9", X"3E", X"03", X"18", X"02", X"3E", X"02", X"CD", --1FC8
  X"30", X"25", X"C4", X"01", X"16", X"CD", X"4D", X"0D", --1FD0
  X"CD", X"DF", X"1F", X"CD", X"EE", X"1B", X"C9", X"DF", --1FD8
  X"CD", X"45", X"20", X"28", X"0D", X"CD", X"4E", X"20", --1FE0
  X"28", X"FB", X"CD", X"FC", X"1F", X"CD", X"4E", X"20", --1FE8
  X"28", X"F3", X"FE", X"29", X"C8", X"CD", X"C3", X"1F", --1FF0
  X"3E", X"0D", X"D7", X"C9", X"DF", X"FE", X"AC", X"20", --1FF8
  X"0D", X"CD", X"79", X"1C", X"CD", X"C3", X"1F", X"CD", --2000
  X"07", X"23", X"3E", X"16", X"18", X"10", X"FE", X"AD", --2008
  X"20", X"12", X"E7", X"CD", X"82", X"1C", X"CD", X"C3", --2010
  X"1F", X"CD", X"99", X"1E", X"3E", X"17", X"D7", X"79", --2018
  X"D7", X"78", X"D7", X"C9", X"CD", X"F2", X"21", X"D0", --2020
  X"CD", X"70", X"20", X"D0", X"CD", X"FB", X"24", X"CD", --2028
  X"C3", X"1F", X"FD", X"CB", X"01", X"76", X"CC", X"F1", --2030
  X"2B", X"C2", X"E3", X"2D", X"78", X"B1", X"0B", X"C8", --2038
  X"1A", X"13", X"D7", X"18", X"F7", X"FE", X"29", X"C8", --2040
  X"FE", X"0D", X"C8", X"FE", X"3A", X"C9", X"DF", X"FE", --2048
  X"3B", X"28", X"14", X"FE", X"2C", X"20", X"0A", X"CD", --2050
  X"30", X"25", X"28", X"0B", X"3E", X"06", X"D7", X"18", --2058
  X"06", X"FE", X"27", X"C0", X"CD", X"F5", X"1F", X"E7", --2060
  X"CD", X"45", X"20", X"20", X"01", X"C1", X"BF", X"C9", --2068
  X"FE", X"23", X"37", X"C0", X"E7", X"CD", X"82", X"1C", --2070
  X"A7", X"CD", X"C3", X"1F", X"CD", X"94", X"1E", X"FE", --2078
  X"10", X"D2", X"0E", X"16", X"CD", X"01", X"16", X"A7", --2080
  X"C9", X"CD", X"30", X"25", X"28", X"08", X"3E", X"01", --2088
  X"CD", X"01", X"16", X"CD", X"6E", X"0D", X"FD", X"36", --2090
  X"02", X"01", X"CD", X"C1", X"20", X"CD", X"EE", X"1B", --2098
  X"ED", X"4B", X"88", X"5C", X"3A", X"6B", X"5C", X"B8", --20A0
  X"38", X"03", X"0E", X"21", X"47", X"ED", X"43", X"88", --20A8
  X"5C", X"3E", X"19", X"90", X"32", X"8C", X"5C", X"FD", --20B0
  X"CB", X"02", X"86", X"CD", X"D9", X"0D", X"C3", X"6E", --20B8
  X"0D", X"CD", X"4E", X"20", X"28", X"FB", X"FE", X"28", --20C0
  X"20", X"0E", X"E7", X"CD", X"DF", X"1F", X"DF", X"FE", --20C8
  X"29", X"C2", X"8A", X"1C", X"E7", X"C3", X"B2", X"21", --20D0
  X"FE", X"CA", X"20", X"11", X"E7", X"CD", X"1F", X"1C", --20D8
  X"FD", X"CB", X"37", X"FE", X"FD", X"CB", X"01", X"76", --20E0
  X"C2", X"8A", X"1C", X"18", X"0D", X"CD", X"8D", X"2C", --20E8
  X"D2", X"AF", X"21", X"CD", X"1F", X"1C", X"FD", X"CB", --20F0
  X"37", X"BE", X"CD", X"30", X"25", X"CA", X"B2", X"21", --20F8
  X"CD", X"BF", X"16", X"21", X"71", X"5C", X"CB", X"B6", --2100
  X"CB", X"EE", X"01", X"01", X"00", X"CB", X"7E", X"20", --2108
  X"0B", X"3A", X"3B", X"5C", X"E6", X"40", X"20", X"02", --2110
  X"0E", X"03", X"B6", X"77", X"F7", X"36", X"0D", X"79", --2118
  X"0F", X"0F", X"30", X"05", X"3E", X"22", X"12", X"2B", --2120
  X"77", X"22", X"5B", X"5C", X"FD", X"CB", X"37", X"7E", --2128
  X"20", X"2C", X"2A", X"5D", X"5C", X"E5", X"2A", X"3D", --2130
  X"5C", X"E5", X"21", X"3A", X"21", X"E5", X"FD", X"CB", --2138
  X"30", X"66", X"28", X"04", X"ED", X"73", X"3D", X"5C", --2140
  X"2A", X"61", X"5C", X"CD", X"A7", X"11", X"FD", X"36", --2148
  X"00", X"FF", X"CD", X"2C", X"0F", X"FD", X"CB", X"01", --2150
  X"BE", X"CD", X"B9", X"21", X"18", X"03", X"CD", X"2C", --2158
  X"0F", X"FD", X"36", X"22", X"00", X"CD", X"D6", X"21", --2160
  X"20", X"0A", X"CD", X"1D", X"11", X"ED", X"4B", X"82", --2168
  X"5C", X"CD", X"D9", X"0D", X"21", X"71", X"5C", X"CB", --2170
  X"AE", X"CB", X"7E", X"CB", X"BE", X"20", X"1C", X"E1", --2178
  X"E1", X"22", X"3D", X"5C", X"E1", X"22", X"5F", X"5C", --2180
  X"FD", X"CB", X"01", X"FE", X"CD", X"B9", X"21", X"2A", --2188
  X"5F", X"5C", X"FD", X"36", X"26", X"00", X"22", X"5D", --2190
  X"5C", X"18", X"17", X"2A", X"63", X"5C", X"ED", X"5B", --2198
  X"61", X"5C", X"37", X"ED", X"52", X"44", X"4D", X"CD", --21A0
  X"B2", X"2A", X"CD", X"FF", X"2A", X"18", X"03", X"CD", --21A8
  X"FC", X"1F", X"CD", X"4E", X"20", X"CA", X"C1", X"20", --21B0
  X"C9", X"2A", X"61", X"5C", X"22", X"5D", X"5C", X"DF", --21B8
  X"FE", X"E2", X"28", X"0C", X"3A", X"71", X"5C", X"CD", --21C0
  X"59", X"1C", X"DF", X"FE", X"0D", X"C8", X"CF", X"0B", --21C8
  X"CD", X"30", X"25", X"C8", X"CF", X"10", X"2A", X"51", --21D0
  X"5C", X"23", X"23", X"23", X"23", X"7E", X"FE", X"4B", --21D8
  X"C9", X"E7", X"CD", X"F2", X"21", X"D8", X"DF", X"FE", --21E0
  X"2C", X"28", X"F6", X"FE", X"3B", X"28", X"F2", X"C3", --21E8
  X"8A", X"1C", X"FE", X"D9", X"D8", X"FE", X"DF", X"3F", --21F0
  X"D8", X"F5", X"E7", X"F1", X"D6", X"C9", X"F5", X"CD", --21F8
  X"82", X"1C", X"F1", X"A7", X"CD", X"C3", X"1F", X"F5", --2200
  X"CD", X"94", X"1E", X"57", X"F1", X"D7", X"7A", X"D7", --2208
  X"C9", X"D6", X"11", X"CE", X"00", X"28", X"1D", X"D6", --2210
  X"02", X"CE", X"00", X"28", X"56", X"FE", X"01", X"7A", --2218
  X"06", X"01", X"20", X"04", X"07", X"07", X"06", X"04", --2220
  X"4F", X"7A", X"FE", X"02", X"30", X"16", X"79", X"21", --2228
  X"91", X"5C", X"18", X"38", X"7A", X"06", X"07", X"38", --2230
  X"05", X"07", X"07", X"07", X"06", X"38", X"4F", X"7A", --2238
  X"FE", X"0A", X"38", X"02", X"CF", X"13", X"21", X"8F", --2240
  X"5C", X"FE", X"08", X"38", X"0B", X"7E", X"28", X"07", --2248
  X"B0", X"2F", X"E6", X"24", X"28", X"01", X"78", X"4F", --2250
  X"79", X"CD", X"6C", X"22", X"3E", X"07", X"BA", X"9F", --2258
  X"CD", X"6C", X"22", X"07", X"07", X"E6", X"50", X"47", --2260
  X"3E", X"08", X"BA", X"9F", X"AE", X"A0", X"AE", X"77", --2268
  X"23", X"78", X"C9", X"9F", X"7A", X"0F", X"06", X"80", --2270
  X"20", X"03", X"0F", X"06", X"40", X"4F", X"7A", X"FE", --2278
  X"08", X"28", X"04", X"FE", X"02", X"30", X"BD", X"79", --2280
  X"21", X"8F", X"5C", X"CD", X"6C", X"22", X"79", X"0F", --2288
  X"0F", X"0F", X"18", X"D8", X"CD", X"94", X"1E", X"FE", --2290
  X"08", X"30", X"A9", X"D3", X"FE", X"07", X"07", X"07", --2298
  X"CB", X"6F", X"20", X"02", X"EE", X"07", X"32", X"48", --22A0
  X"5C", X"C9", X"3E", X"AF", X"90", X"DA", X"F9", X"24", --22A8
  X"47", X"A7", X"1F", X"37", X"1F", X"A7", X"1F", X"A8", --22B0
  X"E6", X"F8", X"A8", X"67", X"79", X"07", X"07", X"07", --22B8
  X"A8", X"E6", X"C7", X"A8", X"07", X"07", X"6F", X"79", --22C0
  X"E6", X"07", X"C9", X"CD", X"07", X"23", X"CD", X"AA", --22C8
  X"22", X"47", X"04", X"7E", X"07", X"10", X"FD", X"E6", --22D0
  X"01", X"C3", X"28", X"2D", X"CD", X"07", X"23", X"CD", --22D8
  X"E5", X"22", X"C3", X"4D", X"0D", X"ED", X"43", X"7D", --22E0
  X"5C", X"CD", X"AA", X"22", X"47", X"04", X"3E", X"FE", --22E8
  X"0F", X"10", X"FD", X"47", X"7E", X"FD", X"4E", X"57", --22F0
  X"CB", X"41", X"20", X"01", X"A0", X"CB", X"51", X"20", --22F8
  X"02", X"A8", X"2F", X"77", X"C3", X"DB", X"0B", X"CD", --2300
  X"14", X"23", X"47", X"C5", X"CD", X"14", X"23", X"59", --2308
  X"C1", X"51", X"4F", X"C9", X"CD", X"D5", X"2D", X"DA", --2310
  X"F9", X"24", X"0E", X"01", X"C8", X"0E", X"FF", X"C9", --2318
  X"DF", X"FE", X"2C", X"C2", X"8A", X"1C", X"E7", X"CD", --2320
  X"82", X"1C", X"CD", X"EE", X"1B", X"EF", X"2A", X"3D", --2328
  X"38", X"7E", X"FE", X"81", X"30", X"05", X"EF", X"02", --2330
  X"38", X"18", X"A1", X"EF", X"A3", X"38", X"36", X"83", --2338
  X"EF", X"C5", X"02", X"38", X"CD", X"7D", X"24", X"C5", --2340
  X"EF", X"31", X"E1", X"04", X"38", X"7E", X"FE", X"80", --2348
  X"30", X"08", X"EF", X"02", X"02", X"38", X"C1", X"C3", --2350
  X"DC", X"22", X"EF", X"C2", X"01", X"C0", X"02", X"03", --2358
  X"01", X"E0", X"0F", X"C0", X"01", X"31", X"E0", X"01", --2360
  X"31", X"E0", X"A0", X"C1", X"02", X"38", X"FD", X"34", --2368
  X"62", X"CD", X"94", X"1E", X"6F", X"E5", X"CD", X"94", --2370
  X"1E", X"E1", X"67", X"22", X"7D", X"5C", X"C1", X"C3", --2378
  X"20", X"24", X"DF", X"FE", X"2C", X"28", X"06", X"CD", --2380
  X"EE", X"1B", X"C3", X"77", X"24", X"E7", X"CD", X"82", --2388
  X"1C", X"CD", X"EE", X"1B", X"EF", X"C5", X"A2", X"04", --2390
  X"1F", X"31", X"30", X"30", X"00", X"06", X"02", X"38", --2398
  X"C3", X"77", X"24", X"C0", X"02", X"C1", X"02", X"31", --23A0
  X"2A", X"E1", X"01", X"E1", X"2A", X"0F", X"E0", X"05", --23A8
  X"2A", X"E0", X"01", X"3D", X"38", X"7E", X"FE", X"81", --23B0
  X"30", X"07", X"EF", X"02", X"02", X"38", X"C3", X"77", --23B8
  X"24", X"CD", X"7D", X"24", X"C5", X"EF", X"02", X"E1", --23C0
  X"01", X"05", X"C1", X"02", X"01", X"31", X"E1", X"04", --23C8
  X"C2", X"02", X"01", X"31", X"E1", X"04", X"E2", X"E5", --23D0
  X"E0", X"03", X"A2", X"04", X"31", X"1F", X"C5", X"02", --23D8
  X"20", X"C0", X"02", X"C2", X"02", X"C1", X"E5", X"04", --23E0
  X"E0", X"E2", X"04", X"0F", X"E1", X"01", X"C1", X"02", --23E8
  X"E0", X"04", X"E2", X"E5", X"04", X"03", X"C2", X"2A", --23F0
  X"E1", X"2A", X"0F", X"02", X"38", X"1A", X"FE", X"81", --23F8
  X"C1", X"DA", X"77", X"24", X"C5", X"EF", X"01", X"38", --2400
  X"3A", X"7D", X"5C", X"CD", X"28", X"2D", X"EF", X"C0", --2408
  X"0F", X"01", X"38", X"3A", X"7E", X"5C", X"CD", X"28", --2410
  X"2D", X"EF", X"C5", X"0F", X"E0", X"E5", X"38", X"C1", --2418
  X"05", X"28", X"3C", X"18", X"14", X"EF", X"E1", X"31", --2420
  X"E3", X"04", X"E2", X"E4", X"04", X"03", X"C1", X"02", --2428
  X"E4", X"04", X"E2", X"E3", X"04", X"0F", X"C2", X"02", --2430
  X"38", X"C5", X"EF", X"C0", X"02", X"E1", X"0F", X"31", --2438
  X"38", X"3A", X"7D", X"5C", X"CD", X"28", X"2D", X"EF", --2440
  X"03", X"E0", X"E2", X"0F", X"C0", X"01", X"E0", X"38", --2448
  X"3A", X"7E", X"5C", X"CD", X"28", X"2D", X"EF", X"03", --2450
  X"38", X"CD", X"B7", X"24", X"C1", X"10", X"C6", X"EF", --2458
  X"02", X"02", X"01", X"38", X"3A", X"7D", X"5C", X"CD", --2460
  X"28", X"2D", X"EF", X"03", X"01", X"38", X"3A", X"7E", --2468
  X"5C", X"CD", X"28", X"2D", X"EF", X"03", X"38", X"CD", --2470
  X"B7", X"24", X"C3", X"4D", X"0D", X"EF", X"31", X"28", --2478
  X"34", X"32", X"00", X"01", X"05", X"E5", X"01", X"05", --2480
  X"2A", X"38", X"CD", X"D5", X"2D", X"38", X"06", X"E6", --2488
  X"FC", X"C6", X"04", X"30", X"02", X"3E", X"FC", X"F5", --2490
  X"CD", X"28", X"2D", X"EF", X"E5", X"01", X"05", X"31", --2498
  X"1F", X"C4", X"02", X"31", X"A2", X"04", X"1F", X"C1", --24A0
  X"01", X"C0", X"02", X"31", X"04", X"31", X"0F", X"A1", --24A8
  X"03", X"1B", X"C3", X"02", X"38", X"C1", X"C9", X"CD", --24B0
  X"07", X"23", X"79", X"B8", X"30", X"06", X"69", X"D5", --24B8
  X"AF", X"5F", X"18", X"07", X"B1", X"C8", X"68", X"41", --24C0
  X"D5", X"16", X"00", X"60", X"78", X"1F", X"85", X"38", --24C8
  X"03", X"BC", X"38", X"07", X"94", X"4F", X"D9", X"C1", --24D0
  X"C5", X"18", X"04", X"4F", X"D5", X"D9", X"C1", X"2A", --24D8
  X"7D", X"5C", X"78", X"84", X"47", X"79", X"3C", X"85", --24E0
  X"38", X"0D", X"28", X"0D", X"3D", X"4F", X"CD", X"E5", --24E8
  X"22", X"D9", X"79", X"10", X"D9", X"D1", X"C9", X"28", --24F0
  X"F3", X"CF", X"0A", X"DF", X"06", X"00", X"C5", X"4F", --24F8
  X"21", X"96", X"25", X"CD", X"DC", X"16", X"79", X"D2", --2500
  X"84", X"26", X"06", X"00", X"4E", X"09", X"E9", X"CD", --2508
  X"74", X"00", X"03", X"FE", X"0D", X"CA", X"8A", X"1C", --2510
  X"FE", X"22", X"20", X"F3", X"CD", X"74", X"00", X"FE", --2518
  X"22", X"C9", X"E7", X"FE", X"28", X"20", X"06", X"CD", --2520
  X"79", X"1C", X"DF", X"FE", X"29", X"C2", X"8A", X"1C", --2528
  X"FD", X"CB", X"01", X"7E", X"C9", X"CD", X"07", X"23", --2530
  X"2A", X"36", X"5C", X"11", X"00", X"01", X"19", X"79", --2538
  X"0F", X"0F", X"0F", X"E6", X"E0", X"A8", X"5F", X"79", --2540
  X"E6", X"18", X"EE", X"40", X"57", X"06", X"60", X"C5", --2548
  X"D5", X"E5", X"1A", X"AE", X"28", X"04", X"3C", X"20", --2550
  X"1A", X"3D", X"4F", X"06", X"07", X"14", X"23", X"1A", --2558
  X"AE", X"A9", X"20", X"0F", X"10", X"F7", X"C1", X"C1", --2560
  X"C1", X"3E", X"80", X"90", X"01", X"01", X"00", X"F7", --2568
  X"12", X"18", X"0A", X"E1", X"11", X"08", X"00", X"19", --2570
  X"D1", X"C1", X"10", X"D3", X"48", X"C3", X"B2", X"2A", --2578
  X"CD", X"07", X"23", X"79", X"0F", X"0F", X"0F", X"4F", --2580
  X"E6", X"E0", X"A8", X"6F", X"79", X"E6", X"03", X"EE", --2588
  X"58", X"67", X"7E", X"C3", X"28", X"2D", X"22", X"1C", --2590
  X"28", X"4F", X"2E", X"F2", X"2B", X"12", X"A8", X"56", --2598
  X"A5", X"57", X"A7", X"84", X"A6", X"8F", X"C4", X"E6", --25A0
  X"AA", X"BF", X"AB", X"C7", X"A9", X"CE", X"00", X"E7", --25A8
  X"C3", X"FF", X"24", X"DF", X"23", X"E5", X"01", X"00", --25B0
  X"00", X"CD", X"0F", X"25", X"20", X"1B", X"CD", X"0F", --25B8
  X"25", X"28", X"FB", X"CD", X"30", X"25", X"28", X"11", --25C0
  X"F7", X"E1", X"D5", X"7E", X"23", X"12", X"13", X"FE", --25C8
  X"22", X"20", X"F8", X"7E", X"23", X"FE", X"22", X"28", --25D0
  X"F2", X"0B", X"D1", X"21", X"3B", X"5C", X"CB", X"B6", --25D8
  X"CB", X"7E", X"C4", X"B2", X"2A", X"C3", X"12", X"27", --25E0
  X"E7", X"CD", X"FB", X"24", X"FE", X"29", X"C2", X"8A", --25E8
  X"1C", X"E7", X"C3", X"12", X"27", X"C3", X"BD", X"27", --25F0
  X"CD", X"30", X"25", X"28", X"28", X"ED", X"4B", X"76", --25F8
  X"5C", X"CD", X"2B", X"2D", X"EF", X"A1", X"0F", X"34", --2600
  X"37", X"16", X"04", X"34", X"80", X"41", X"00", X"00", --2608
  X"80", X"32", X"02", X"A1", X"03", X"31", X"38", X"CD", --2610
  X"A2", X"2D", X"ED", X"43", X"76", X"5C", X"7E", X"A7", --2618
  X"28", X"03", X"D6", X"10", X"77", X"18", X"09", X"CD", --2620
  X"30", X"25", X"28", X"04", X"EF", X"A3", X"38", X"34", --2628
  X"E7", X"C3", X"C3", X"26", X"01", X"5A", X"10", X"E7", --2630
  X"FE", X"23", X"CA", X"0D", X"27", X"21", X"3B", X"5C", --2638
  X"CB", X"B6", X"CB", X"7E", X"28", X"1F", X"CD", X"8E", --2640
  X"02", X"0E", X"00", X"20", X"13", X"CD", X"1E", X"03", --2648
  X"30", X"0E", X"15", X"5F", X"CD", X"33", X"03", X"F5", --2650
  X"01", X"01", X"00", X"F7", X"F1", X"12", X"0E", X"01", --2658
  X"06", X"00", X"CD", X"B2", X"2A", X"C3", X"12", X"27", --2660
  X"CD", X"22", X"25", X"C4", X"35", X"25", X"E7", X"C3", --2668
  X"DB", X"25", X"CD", X"22", X"25", X"C4", X"80", X"25", --2670
  X"E7", X"18", X"48", X"CD", X"22", X"25", X"C4", X"CB", --2678
  X"22", X"E7", X"18", X"3F", X"CD", X"88", X"2C", X"30", --2680
  X"56", X"FE", X"41", X"30", X"3C", X"CD", X"30", X"25", --2688
  X"20", X"23", X"CD", X"9B", X"2C", X"DF", X"01", X"06", --2690
  X"00", X"CD", X"55", X"16", X"23", X"36", X"0E", X"23", --2698
  X"EB", X"2A", X"65", X"5C", X"0E", X"05", X"A7", X"ED", --26A0
  X"42", X"22", X"65", X"5C", X"ED", X"B0", X"EB", X"2B", --26A8
  X"CD", X"77", X"00", X"18", X"0E", X"DF", X"23", X"7E", --26B0
  X"FE", X"0E", X"20", X"FA", X"23", X"CD", X"B4", X"33", --26B8
  X"22", X"5D", X"5C", X"FD", X"CB", X"01", X"F6", X"18", --26C0
  X"14", X"CD", X"B2", X"28", X"DA", X"2E", X"1C", X"CC", --26C8
  X"96", X"29", X"3A", X"3B", X"5C", X"FE", X"C0", X"38", --26D0
  X"04", X"23", X"CD", X"B4", X"33", X"18", X"33", X"01", --26D8
  X"DB", X"09", X"FE", X"2D", X"28", X"27", X"01", X"18", --26E0
  X"10", X"FE", X"AE", X"28", X"20", X"D6", X"AF", X"DA", --26E8
  X"8A", X"1C", X"01", X"F0", X"04", X"FE", X"14", X"28", --26F0
  X"14", X"D2", X"8A", X"1C", X"06", X"10", X"C6", X"DC", --26F8
  X"4F", X"FE", X"DF", X"30", X"02", X"CB", X"B1", X"FE", --2700
  X"EE", X"38", X"02", X"CB", X"B9", X"C5", X"E7", X"C3", --2708
  X"FF", X"24", X"DF", X"FE", X"28", X"20", X"0C", X"FD", --2710
  X"CB", X"01", X"76", X"20", X"17", X"CD", X"52", X"2A", --2718
  X"E7", X"18", X"F0", X"06", X"00", X"4F", X"21", X"95", --2720
  X"27", X"CD", X"DC", X"16", X"30", X"06", X"4E", X"21", --2728
  X"ED", X"26", X"09", X"46", X"D1", X"7A", X"B8", X"38", --2730
  X"3A", X"A7", X"CA", X"18", X"00", X"C5", X"21", X"3B", --2738
  X"5C", X"7B", X"FE", X"ED", X"20", X"06", X"CB", X"76", --2740
  X"20", X"02", X"1E", X"99", X"D5", X"CD", X"30", X"25", --2748
  X"28", X"09", X"7B", X"E6", X"3F", X"47", X"EF", X"3B", --2750
  X"38", X"18", X"09", X"7B", X"FD", X"AE", X"01", X"E6", --2758
  X"40", X"C2", X"8A", X"1C", X"D1", X"21", X"3B", X"5C", --2760
  X"CB", X"F6", X"CB", X"7B", X"20", X"02", X"CB", X"B6", --2768
  X"C1", X"18", X"C1", X"D5", X"79", X"FD", X"CB", X"01", --2770
  X"76", X"20", X"15", X"E6", X"3F", X"C6", X"08", X"4F", --2778
  X"FE", X"10", X"20", X"04", X"CB", X"F1", X"18", X"08", --2780
  X"38", X"D7", X"FE", X"17", X"28", X"02", X"CB", X"F9", --2788
  X"C5", X"E7", X"C3", X"FF", X"24", X"2B", X"CF", X"2D", --2790
  X"C3", X"2A", X"C4", X"2F", X"C5", X"5E", X"C6", X"3D", --2798
  X"CE", X"3E", X"CC", X"3C", X"CD", X"C7", X"C9", X"C8", --27A0
  X"CA", X"C9", X"CB", X"C5", X"C7", X"C6", X"C8", X"00", --27A8
  X"06", X"08", X"08", X"0A", X"02", X"03", X"05", X"05", --27B0
  X"05", X"05", X"05", X"05", X"06", X"CD", X"30", X"25", --27B8
  X"20", X"35", X"E7", X"CD", X"8D", X"2C", X"D2", X"8A", --27C0
  X"1C", X"E7", X"FE", X"24", X"F5", X"20", X"01", X"E7", --27C8
  X"FE", X"28", X"20", X"12", X"E7", X"FE", X"29", X"28", --27D0
  X"10", X"CD", X"FB", X"24", X"DF", X"FE", X"2C", X"20", --27D8
  X"03", X"E7", X"18", X"F5", X"FE", X"29", X"C2", X"8A", --27E0
  X"1C", X"E7", X"21", X"3B", X"5C", X"CB", X"B6", X"F1", --27E8
  X"28", X"02", X"CB", X"F6", X"C3", X"12", X"27", X"E7", --27F0
  X"E6", X"DF", X"47", X"E7", X"D6", X"24", X"4F", X"20", --27F8
  X"01", X"E7", X"E7", X"E5", X"2A", X"53", X"5C", X"2B", --2800
  X"11", X"CE", X"00", X"C5", X"CD", X"86", X"1D", X"C1", --2808
  X"30", X"02", X"CF", X"18", X"E5", X"CD", X"AB", X"28", --2810
  X"E6", X"DF", X"B8", X"20", X"08", X"CD", X"AB", X"28", --2818
  X"D6", X"24", X"B9", X"28", X"0C", X"E1", X"2B", X"11", --2820
  X"00", X"02", X"C5", X"CD", X"8B", X"19", X"C1", X"18", --2828
  X"D7", X"A7", X"CC", X"AB", X"28", X"D1", X"D1", X"ED", --2830
  X"53", X"5D", X"5C", X"CD", X"AB", X"28", X"E5", X"FE", --2838
  X"29", X"28", X"42", X"23", X"7E", X"FE", X"0E", X"16", --2840
  X"40", X"28", X"07", X"2B", X"CD", X"AB", X"28", X"23", --2848
  X"16", X"00", X"23", X"E5", X"D5", X"CD", X"FB", X"24", --2850
  X"F1", X"FD", X"AE", X"01", X"E6", X"40", X"20", X"2B", --2858
  X"E1", X"EB", X"2A", X"65", X"5C", X"01", X"05", X"00", --2860
  X"ED", X"42", X"22", X"65", X"5C", X"ED", X"B0", X"EB", --2868
  X"2B", X"CD", X"AB", X"28", X"FE", X"29", X"28", X"0D", --2870
  X"E5", X"DF", X"FE", X"2C", X"20", X"0D", X"E7", X"E1", --2878
  X"CD", X"AB", X"28", X"18", X"BE", X"E5", X"DF", X"FE", --2880
  X"29", X"28", X"02", X"CF", X"19", X"D1", X"EB", X"22", --2888
  X"5D", X"5C", X"2A", X"0B", X"5C", X"E3", X"22", X"0B", --2890
  X"5C", X"D5", X"E7", X"E7", X"CD", X"FB", X"24", X"E1", --2898
  X"22", X"5D", X"5C", X"E1", X"22", X"0B", X"5C", X"E7", --28A0
  X"C3", X"12", X"27", X"23", X"7E", X"FE", X"21", X"38", --28A8
  X"FA", X"C9", X"FD", X"CB", X"01", X"F6", X"DF", X"CD", --28B0
  X"8D", X"2C", X"D2", X"8A", X"1C", X"E5", X"E6", X"1F", --28B8
  X"4F", X"E7", X"E5", X"FE", X"28", X"28", X"28", X"CB", --28C0
  X"F1", X"FE", X"24", X"28", X"11", X"CB", X"E9", X"CD", --28C8
  X"88", X"2C", X"30", X"0F", X"CD", X"88", X"2C", X"30", --28D0
  X"16", X"CB", X"B1", X"E7", X"18", X"F6", X"E7", X"FD", --28D8
  X"CB", X"01", X"B6", X"3A", X"0C", X"5C", X"A7", X"28", --28E0
  X"06", X"CD", X"30", X"25", X"C2", X"51", X"29", X"41", --28E8
  X"CD", X"30", X"25", X"20", X"08", X"79", X"E6", X"E0", --28F0
  X"CB", X"FF", X"4F", X"18", X"37", X"2A", X"4B", X"5C", --28F8
  X"7E", X"E6", X"7F", X"28", X"2D", X"B9", X"20", X"22", --2900
  X"17", X"87", X"F2", X"3F", X"29", X"38", X"30", X"D1", --2908
  X"D5", X"E5", X"23", X"1A", X"13", X"FE", X"20", X"28", --2910
  X"FA", X"F6", X"20", X"BE", X"28", X"F4", X"F6", X"80", --2918
  X"BE", X"20", X"06", X"1A", X"CD", X"88", X"2C", X"30", --2920
  X"15", X"E1", X"C5", X"CD", X"B8", X"19", X"EB", X"C1", --2928
  X"18", X"CE", X"CB", X"F8", X"D1", X"DF", X"FE", X"28", --2930
  X"28", X"09", X"CB", X"E8", X"18", X"0D", X"D1", X"D1", --2938
  X"D1", X"E5", X"DF", X"CD", X"88", X"2C", X"30", X"03", --2940
  X"E7", X"18", X"F8", X"E1", X"CB", X"10", X"CB", X"70", --2948
  X"C9", X"2A", X"0B", X"5C", X"7E", X"FE", X"29", X"CA", --2950
  X"EF", X"28", X"7E", X"F6", X"60", X"47", X"23", X"7E", --2958
  X"FE", X"0E", X"28", X"07", X"2B", X"CD", X"AB", X"28", --2960
  X"23", X"CB", X"A8", X"78", X"B9", X"28", X"12", X"23", --2968
  X"23", X"23", X"23", X"23", X"CD", X"AB", X"28", X"FE", --2970
  X"29", X"CA", X"EF", X"28", X"CD", X"AB", X"28", X"18", --2978
  X"D9", X"CB", X"69", X"20", X"0C", X"23", X"ED", X"5B", --2980
  X"65", X"5C", X"CD", X"C0", X"33", X"EB", X"22", X"65", --2988
  X"5C", X"D1", X"D1", X"AF", X"3C", X"C9", X"AF", X"47", --2990
  X"CB", X"79", X"20", X"4B", X"CB", X"7E", X"20", X"0E", --2998
  X"3C", X"23", X"4E", X"23", X"46", X"23", X"EB", X"CD", --29A0
  X"B2", X"2A", X"DF", X"C3", X"49", X"2A", X"23", X"23", --29A8
  X"23", X"46", X"CB", X"71", X"28", X"0A", X"05", X"28", --29B0
  X"E8", X"EB", X"DF", X"FE", X"28", X"20", X"61", X"EB", --29B8
  X"EB", X"18", X"24", X"E5", X"DF", X"E1", X"FE", X"2C", --29C0
  X"28", X"20", X"CB", X"79", X"28", X"52", X"CB", X"71", --29C8
  X"20", X"06", X"FE", X"29", X"20", X"3C", X"E7", X"C9", --29D0
  X"FE", X"29", X"28", X"6C", X"FE", X"CC", X"20", X"32", --29D8
  X"DF", X"2B", X"22", X"5D", X"5C", X"18", X"5E", X"21", --29E0
  X"00", X"00", X"E5", X"E7", X"E1", X"79", X"FE", X"C0", --29E8
  X"20", X"09", X"DF", X"FE", X"29", X"28", X"51", X"FE", --29F0
  X"CC", X"28", X"E5", X"C5", X"E5", X"CD", X"EE", X"2A", --29F8
  X"E3", X"EB", X"CD", X"CC", X"2A", X"38", X"19", X"0B", --2A00
  X"CD", X"F4", X"2A", X"09", X"D1", X"C1", X"10", X"B3", --2A08
  X"CB", X"79", X"20", X"66", X"E5", X"CB", X"71", X"20", --2A10
  X"13", X"42", X"4B", X"DF", X"FE", X"29", X"28", X"02", --2A18
  X"CF", X"02", X"E7", X"E1", X"11", X"05", X"00", X"CD", --2A20
  X"F4", X"2A", X"09", X"C9", X"CD", X"EE", X"2A", X"E3", --2A28
  X"CD", X"F4", X"2A", X"C1", X"09", X"23", X"42", X"4B", --2A30
  X"EB", X"CD", X"B1", X"2A", X"DF", X"FE", X"29", X"28", --2A38
  X"07", X"FE", X"2C", X"20", X"DB", X"CD", X"52", X"2A", --2A40
  X"E7", X"FE", X"28", X"28", X"F8", X"FD", X"CB", X"01", --2A48
  X"B6", X"C9", X"CD", X"30", X"25", X"C4", X"F1", X"2B", --2A50
  X"E7", X"FE", X"29", X"28", X"50", X"D5", X"AF", X"F5", --2A58
  X"C5", X"11", X"01", X"00", X"DF", X"E1", X"FE", X"CC", --2A60
  X"28", X"17", X"F1", X"CD", X"CD", X"2A", X"F5", X"50", --2A68
  X"59", X"E5", X"DF", X"E1", X"FE", X"CC", X"28", X"09", --2A70
  X"FE", X"29", X"C2", X"8A", X"1C", X"62", X"6B", X"18", --2A78
  X"13", X"E5", X"E7", X"E1", X"FE", X"29", X"28", X"0C", --2A80
  X"F1", X"CD", X"CD", X"2A", X"F5", X"DF", X"60", X"69", --2A88
  X"FE", X"29", X"20", X"E6", X"F1", X"E3", X"19", X"2B", --2A90
  X"E3", X"A7", X"ED", X"52", X"01", X"00", X"00", X"38", --2A98
  X"07", X"23", X"A7", X"FA", X"20", X"2A", X"44", X"4D", --2AA0
  X"D1", X"FD", X"CB", X"01", X"B6", X"CD", X"30", X"25", --2AA8
  X"C8", X"AF", X"FD", X"CB", X"01", X"B6", X"C5", X"CD", --2AB0
  X"A9", X"33", X"C1", X"2A", X"65", X"5C", X"77", X"23", --2AB8
  X"73", X"23", X"72", X"23", X"71", X"23", X"70", X"23", --2AC0
  X"22", X"65", X"5C", X"C9", X"AF", X"D5", X"E5", X"F5", --2AC8
  X"CD", X"82", X"1C", X"F1", X"CD", X"30", X"25", X"28", --2AD0
  X"12", X"F5", X"CD", X"99", X"1E", X"D1", X"78", X"B1", --2AD8
  X"37", X"28", X"05", X"E1", X"E5", X"A7", X"ED", X"42", --2AE0
  X"7A", X"DE", X"00", X"E1", X"D1", X"C9", X"EB", X"23", --2AE8
  X"5E", X"23", X"56", X"C9", X"CD", X"30", X"25", X"C8", --2AF0
  X"CD", X"A9", X"30", X"DA", X"15", X"1F", X"C9", X"2A", --2AF8
  X"4D", X"5C", X"FD", X"CB", X"37", X"4E", X"28", X"5E", --2B00
  X"01", X"05", X"00", X"03", X"23", X"7E", X"FE", X"20", --2B08
  X"28", X"FA", X"30", X"0B", X"FE", X"10", X"38", X"11", --2B10
  X"FE", X"16", X"30", X"0D", X"23", X"18", X"ED", X"CD", --2B18
  X"88", X"2C", X"38", X"E7", X"FE", X"24", X"CA", X"C0", --2B20
  X"2B", X"79", X"2A", X"59", X"5C", X"2B", X"CD", X"55", --2B28
  X"16", X"23", X"23", X"EB", X"D5", X"2A", X"4D", X"5C", --2B30
  X"1B", X"D6", X"06", X"47", X"28", X"11", X"23", X"7E", --2B38
  X"FE", X"21", X"38", X"FA", X"F6", X"20", X"13", X"12", --2B40
  X"10", X"F4", X"F6", X"80", X"12", X"3E", X"C0", X"2A", --2B48
  X"4D", X"5C", X"AE", X"F6", X"20", X"E1", X"CD", X"EA", --2B50
  X"2B", X"E5", X"EF", X"02", X"38", X"E1", X"01", X"05", --2B58
  X"00", X"A7", X"ED", X"42", X"18", X"40", X"FD", X"CB", --2B60
  X"01", X"76", X"28", X"06", X"11", X"06", X"00", X"19", --2B68
  X"18", X"E7", X"2A", X"4D", X"5C", X"ED", X"4B", X"72", --2B70
  X"5C", X"FD", X"CB", X"37", X"46", X"20", X"30", X"78", --2B78
  X"B1", X"C8", X"E5", X"F7", X"D5", X"C5", X"54", X"5D", --2B80
  X"23", X"36", X"20", X"ED", X"B8", X"E5", X"CD", X"F1", --2B88
  X"2B", X"E1", X"E3", X"A7", X"ED", X"42", X"09", X"30", --2B90
  X"02", X"44", X"4D", X"E3", X"EB", X"78", X"B1", X"28", --2B98
  X"02", X"ED", X"B0", X"C1", X"D1", X"E1", X"EB", X"78", --2BA0
  X"B1", X"C8", X"D5", X"ED", X"B0", X"E1", X"C9", X"2B", --2BA8
  X"2B", X"2B", X"7E", X"E5", X"C5", X"CD", X"C6", X"2B", --2BB0
  X"C1", X"E1", X"03", X"03", X"03", X"C3", X"E8", X"19", --2BB8
  X"3E", X"DF", X"2A", X"4D", X"5C", X"A6", X"F5", X"CD", --2BC0
  X"F1", X"2B", X"EB", X"09", X"C5", X"2B", X"22", X"4D", --2BC8
  X"5C", X"03", X"03", X"03", X"2A", X"59", X"5C", X"2B", --2BD0
  X"CD", X"55", X"16", X"2A", X"4D", X"5C", X"C1", X"C5", --2BD8
  X"03", X"ED", X"B8", X"EB", X"23", X"C1", X"70", X"2B", --2BE0
  X"71", X"F1", X"2B", X"77", X"2A", X"59", X"5C", X"2B", --2BE8
  X"C9", X"2A", X"65", X"5C", X"2B", X"46", X"2B", X"4E", --2BF0
  X"2B", X"56", X"2B", X"5E", X"2B", X"7E", X"22", X"65", --2BF8
  X"5C", X"C9", X"CD", X"B2", X"28", X"C2", X"8A", X"1C", --2C00
  X"CD", X"30", X"25", X"20", X"08", X"CB", X"B1", X"CD", --2C08
  X"96", X"29", X"CD", X"EE", X"1B", X"38", X"08", X"C5", --2C10
  X"CD", X"B8", X"19", X"CD", X"E8", X"19", X"C1", X"CB", --2C18
  X"F9", X"06", X"00", X"C5", X"21", X"01", X"00", X"CB", --2C20
  X"71", X"20", X"02", X"2E", X"05", X"EB", X"E7", X"26", --2C28
  X"FF", X"CD", X"CC", X"2A", X"DA", X"20", X"2A", X"E1", --2C30
  X"C5", X"24", X"E5", X"60", X"69", X"CD", X"F4", X"2A", --2C38
  X"EB", X"DF", X"FE", X"2C", X"28", X"E8", X"FE", X"29", --2C40
  X"20", X"BB", X"E7", X"C1", X"79", X"68", X"26", X"00", --2C48
  X"23", X"23", X"29", X"19", X"DA", X"15", X"1F", X"D5", --2C50
  X"C5", X"E5", X"44", X"4D", X"2A", X"59", X"5C", X"2B", --2C58
  X"CD", X"55", X"16", X"23", X"77", X"C1", X"0B", X"0B", --2C60
  X"0B", X"23", X"71", X"23", X"70", X"C1", X"78", X"23", --2C68
  X"77", X"62", X"6B", X"1B", X"36", X"00", X"CB", X"71", --2C70
  X"28", X"02", X"36", X"20", X"C1", X"ED", X"B8", X"C1", --2C78
  X"70", X"2B", X"71", X"2B", X"3D", X"20", X"F8", X"C9", --2C80
  X"CD", X"1B", X"2D", X"3F", X"D8", X"FE", X"41", X"3F", --2C88
  X"D0", X"FE", X"5B", X"D8", X"FE", X"61", X"3F", X"D0", --2C90
  X"FE", X"7B", X"C9", X"FE", X"C4", X"20", X"19", X"11", --2C98
  X"00", X"00", X"E7", X"D6", X"31", X"CE", X"00", X"20", --2CA0
  X"0A", X"EB", X"3F", X"ED", X"6A", X"DA", X"AD", X"31", --2CA8
  X"EB", X"18", X"EF", X"42", X"4B", X"C3", X"2B", X"2D", --2CB0
  X"FE", X"2E", X"28", X"0F", X"CD", X"3B", X"2D", X"FE", --2CB8
  X"2E", X"20", X"28", X"E7", X"CD", X"1B", X"2D", X"38", --2CC0
  X"22", X"18", X"0A", X"E7", X"CD", X"1B", X"2D", X"DA", --2CC8
  X"8A", X"1C", X"EF", X"A0", X"38", X"EF", X"A1", X"C0", --2CD0
  X"02", X"38", X"DF", X"CD", X"22", X"2D", X"38", X"0B", --2CD8
  X"EF", X"E0", X"A4", X"05", X"C0", X"04", X"0F", X"38", --2CE0
  X"E7", X"18", X"EF", X"FE", X"45", X"28", X"03", X"FE", --2CE8
  X"65", X"C0", X"06", X"FF", X"E7", X"FE", X"2B", X"28", --2CF0
  X"05", X"FE", X"2D", X"20", X"02", X"04", X"E7", X"CD", --2CF8
  X"1B", X"2D", X"38", X"CB", X"C5", X"CD", X"3B", X"2D", --2D00
  X"CD", X"D5", X"2D", X"C1", X"DA", X"AD", X"31", X"A7", --2D08
  X"FA", X"AD", X"31", X"04", X"28", X"02", X"ED", X"44", --2D10
  X"C3", X"4F", X"2D", X"FE", X"30", X"D8", X"FE", X"3A", --2D18
  X"3F", X"C9", X"CD", X"1B", X"2D", X"D8", X"D6", X"30", --2D20
  X"4F", X"06", X"00", X"FD", X"21", X"3A", X"5C", X"AF", --2D28
  X"5F", X"51", X"48", X"47", X"CD", X"B6", X"2A", X"EF", --2D30
  X"38", X"A7", X"C9", X"F5", X"EF", X"A0", X"38", X"F1", --2D38
  X"CD", X"22", X"2D", X"D8", X"EF", X"01", X"A4", X"04", --2D40
  X"0F", X"38", X"CD", X"74", X"00", X"18", X"F1", X"07", --2D48
  X"0F", X"30", X"02", X"2F", X"3C", X"F5", X"21", X"92", --2D50
  X"5C", X"CD", X"0B", X"35", X"EF", X"A4", X"38", X"F1", --2D58
  X"CB", X"3F", X"30", X"0D", X"F5", X"EF", X"C1", X"E0", --2D60
  X"00", X"04", X"04", X"33", X"02", X"05", X"E1", X"38", --2D68
  X"F1", X"28", X"08", X"F5", X"EF", X"31", X"04", X"38", --2D70
  X"F1", X"18", X"E5", X"EF", X"02", X"38", X"C9", X"23", --2D78
  X"4E", X"23", X"7E", X"A9", X"91", X"5F", X"23", X"7E", --2D80
  X"89", X"A9", X"57", X"C9", X"0E", X"00", X"E5", X"36", --2D88
  X"00", X"23", X"71", X"23", X"7B", X"A9", X"91", X"77", --2D90
  X"23", X"7A", X"89", X"A9", X"77", X"23", X"36", X"00", --2D98
  X"E1", X"C9", X"EF", X"38", X"7E", X"A7", X"28", X"05", --2DA0
  X"EF", X"A2", X"0F", X"27", X"38", X"EF", X"02", X"38", --2DA8
  X"E5", X"D5", X"EB", X"46", X"CD", X"7F", X"2D", X"AF", --2DB0
  X"90", X"CB", X"79", X"42", X"4B", X"7B", X"D1", X"E1", --2DB8
  X"C9", X"57", X"17", X"9F", X"5F", X"4F", X"AF", X"47", --2DC0
  X"CD", X"B6", X"2A", X"EF", X"34", X"EF", X"1A", X"20", --2DC8
  X"9A", X"85", X"04", X"27", X"38", X"CD", X"A2", X"2D", --2DD0
  X"D8", X"F5", X"05", X"04", X"28", X"03", X"F1", X"37", --2DD8
  X"C9", X"F1", X"C9", X"EF", X"31", X"36", X"00", X"0B", --2DE0
  X"31", X"37", X"00", X"0D", X"02", X"38", X"3E", X"30", --2DE8
  X"D7", X"C9", X"2A", X"38", X"3E", X"2D", X"D7", X"EF", --2DF0
  X"A0", X"C3", X"C4", X"C5", X"02", X"38", X"D9", X"E5", --2DF8
  X"D9", X"EF", X"31", X"27", X"C2", X"03", X"E2", X"01", --2E00
  X"C2", X"02", X"38", X"7E", X"A7", X"20", X"47", X"CD", --2E08
  X"7F", X"2D", X"06", X"10", X"7A", X"A7", X"20", X"06", --2E10
  X"B3", X"28", X"09", X"53", X"06", X"08", X"D5", X"D9", --2E18
  X"D1", X"D9", X"18", X"57", X"EF", X"E2", X"38", X"7E", --2E20
  X"D6", X"7E", X"CD", X"C1", X"2D", X"57", X"3A", X"AC", --2E28
  X"5C", X"92", X"32", X"AC", X"5C", X"7A", X"CD", X"4F", --2E30
  X"2D", X"EF", X"31", X"27", X"C1", X"03", X"E1", X"38", --2E38
  X"CD", X"D5", X"2D", X"E5", X"32", X"A1", X"5C", X"3D", --2E40
  X"17", X"9F", X"3C", X"21", X"AB", X"5C", X"77", X"23", --2E48
  X"86", X"77", X"E1", X"C3", X"CF", X"2E", X"D6", X"80", --2E50
  X"FE", X"1C", X"38", X"13", X"CD", X"C1", X"2D", X"D6", --2E58
  X"07", X"47", X"21", X"AC", X"5C", X"86", X"77", X"78", --2E60
  X"ED", X"44", X"CD", X"4F", X"2D", X"18", X"92", X"EB", --2E68
  X"CD", X"BA", X"2F", X"D9", X"CB", X"FA", X"7D", X"D9", --2E70
  X"D6", X"80", X"47", X"CB", X"23", X"CB", X"12", X"D9", --2E78
  X"CB", X"13", X"CB", X"12", X"D9", X"21", X"AA", X"5C", --2E80
  X"0E", X"05", X"7E", X"8F", X"27", X"77", X"2B", X"0D", --2E88
  X"20", X"F8", X"10", X"E7", X"AF", X"21", X"A6", X"5C", --2E90
  X"11", X"A1", X"5C", X"06", X"09", X"ED", X"6F", X"0E", --2E98
  X"FF", X"ED", X"6F", X"20", X"04", X"0D", X"0C", X"20", --2EA0
  X"0A", X"12", X"13", X"FD", X"34", X"71", X"FD", X"34", --2EA8
  X"72", X"0E", X"00", X"CB", X"40", X"28", X"01", X"23", --2EB0
  X"10", X"E7", X"3A", X"AB", X"5C", X"D6", X"09", X"38", --2EB8
  X"0A", X"FD", X"35", X"71", X"3E", X"04", X"FD", X"BE", --2EC0
  X"6F", X"18", X"41", X"EF", X"02", X"E2", X"38", X"EB", --2EC8
  X"CD", X"BA", X"2F", X"D9", X"3E", X"80", X"95", X"2E", --2ED0
  X"00", X"CB", X"FA", X"D9", X"CD", X"DD", X"2F", X"FD", --2ED8
  X"7E", X"71", X"FE", X"08", X"38", X"06", X"D9", X"CB", --2EE0
  X"12", X"D9", X"18", X"20", X"01", X"00", X"02", X"7B", --2EE8
  X"CD", X"8B", X"2F", X"5F", X"7A", X"CD", X"8B", X"2F", --2EF0
  X"57", X"C5", X"D9", X"C1", X"10", X"F1", X"21", X"A1", --2EF8
  X"5C", X"79", X"FD", X"4E", X"71", X"09", X"77", X"FD", --2F00
  X"34", X"71", X"18", X"D3", X"F5", X"21", X"A1", X"5C", --2F08
  X"FD", X"4E", X"71", X"06", X"00", X"09", X"41", X"F1", --2F10
  X"2B", X"7E", X"CE", X"00", X"77", X"A7", X"28", X"05", --2F18
  X"FE", X"0A", X"3F", X"30", X"08", X"10", X"F1", X"36", --2F20
  X"01", X"04", X"FD", X"34", X"72", X"FD", X"70", X"71", --2F28
  X"EF", X"02", X"38", X"D9", X"E1", X"D9", X"ED", X"4B", --2F30
  X"AB", X"5C", X"21", X"A1", X"5C", X"78", X"FE", X"09", --2F38
  X"38", X"04", X"FE", X"FC", X"38", X"26", X"A7", X"CC", --2F40
  X"EF", X"15", X"AF", X"90", X"FA", X"52", X"2F", X"47", --2F48
  X"18", X"0C", X"79", X"A7", X"28", X"03", X"7E", X"23", --2F50
  X"0D", X"CD", X"EF", X"15", X"10", X"F4", X"79", X"A7", --2F58
  X"C8", X"04", X"3E", X"2E", X"D7", X"3E", X"30", X"10", --2F60
  X"FB", X"41", X"18", X"E6", X"50", X"15", X"06", X"01", --2F68
  X"CD", X"4A", X"2F", X"3E", X"45", X"D7", X"4A", X"79", --2F70
  X"A7", X"F2", X"83", X"2F", X"ED", X"44", X"4F", X"3E", --2F78
  X"2D", X"18", X"02", X"3E", X"2B", X"D7", X"06", X"00", --2F80
  X"C3", X"1B", X"1A", X"D5", X"6F", X"26", X"00", X"5D", --2F88
  X"54", X"29", X"29", X"19", X"29", X"59", X"19", X"4C", --2F90
  X"7D", X"D1", X"C9", X"7E", X"36", X"00", X"A7", X"C8", --2F98
  X"23", X"CB", X"7E", X"CB", X"FE", X"2B", X"C8", X"C5", --2FA0
  X"01", X"05", X"00", X"09", X"41", X"4F", X"37", X"2B", --2FA8
  X"7E", X"2F", X"CE", X"00", X"77", X"10", X"F8", X"79", --2FB0
  X"C1", X"C9", X"E5", X"F5", X"4E", X"23", X"46", X"77", --2FB8
  X"23", X"79", X"4E", X"C5", X"23", X"4E", X"23", X"46", --2FC0
  X"EB", X"57", X"5E", X"D5", X"23", X"56", X"23", X"5E", --2FC8
  X"D5", X"D9", X"D1", X"E1", X"C1", X"D9", X"23", X"56", --2FD0
  X"23", X"5E", X"F1", X"E1", X"C9", X"A7", X"C8", X"FE", --2FD8
  X"21", X"30", X"16", X"C5", X"47", X"D9", X"CB", X"2D", --2FE0
  X"CB", X"1A", X"CB", X"1B", X"D9", X"CB", X"1A", X"CB", --2FE8
  X"1B", X"10", X"F2", X"C1", X"D0", X"CD", X"04", X"30", --2FF0
  X"C0", X"D9", X"AF", X"2E", X"00", X"57", X"5D", X"D9", --2FF8
  X"11", X"00", X"00", X"C9", X"1C", X"C0", X"14", X"C0", --3000
  X"D9", X"1C", X"20", X"01", X"14", X"D9", X"C9", X"EB", --3008
  X"CD", X"6E", X"34", X"EB", X"1A", X"B6", X"20", X"26", --3010
  X"D5", X"23", X"E5", X"23", X"5E", X"23", X"56", X"23", --3018
  X"23", X"23", X"7E", X"23", X"4E", X"23", X"46", X"E1", --3020
  X"EB", X"09", X"EB", X"8E", X"0F", X"CE", X"00", X"20", --3028
  X"0B", X"9F", X"77", X"23", X"73", X"23", X"72", X"2B", --3030
  X"2B", X"2B", X"D1", X"C9", X"2B", X"D1", X"CD", X"93", --3038
  X"32", X"D9", X"E5", X"D9", X"D5", X"E5", X"CD", X"9B", --3040
  X"2F", X"47", X"EB", X"CD", X"9B", X"2F", X"4F", X"B8", --3048
  X"30", X"03", X"78", X"41", X"EB", X"F5", X"90", X"CD", --3050
  X"BA", X"2F", X"CD", X"DD", X"2F", X"F1", X"E1", X"77", --3058
  X"E5", X"68", X"61", X"19", X"D9", X"EB", X"ED", X"4A", --3060
  X"EB", X"7C", X"8D", X"6F", X"1F", X"AD", X"D9", X"EB", --3068
  X"E1", X"1F", X"30", X"08", X"3E", X"01", X"CD", X"DD", --3070
  X"2F", X"34", X"28", X"23", X"D9", X"7D", X"E6", X"80", --3078
  X"D9", X"23", X"77", X"2B", X"28", X"1F", X"7B", X"ED", --3080
  X"44", X"3F", X"5F", X"7A", X"2F", X"CE", X"00", X"57", --3088
  X"D9", X"7B", X"2F", X"CE", X"00", X"5F", X"7A", X"2F", --3090
  X"CE", X"00", X"30", X"07", X"1F", X"D9", X"34", X"CA", --3098
  X"AD", X"31", X"D9", X"57", X"D9", X"AF", X"C3", X"55", --30A0
  X"31", X"C5", X"06", X"10", X"7C", X"4D", X"21", X"00", --30A8
  X"00", X"29", X"38", X"0A", X"CB", X"11", X"17", X"30", --30B0
  X"03", X"19", X"38", X"02", X"10", X"F3", X"C1", X"C9", --30B8
  X"CD", X"E9", X"34", X"D8", X"23", X"AE", X"CB", X"FE", --30C0
  X"2B", X"C9", X"1A", X"B6", X"20", X"22", X"D5", X"E5", --30C8
  X"D5", X"CD", X"7F", X"2D", X"EB", X"E3", X"41", X"CD", --30D0
  X"7F", X"2D", X"78", X"A9", X"4F", X"E1", X"CD", X"A9", --30D8
  X"30", X"EB", X"E1", X"38", X"0A", X"7A", X"B3", X"20", --30E0
  X"01", X"4F", X"CD", X"8E", X"2D", X"D1", X"C9", X"D1", --30E8
  X"CD", X"93", X"32", X"AF", X"CD", X"C0", X"30", X"D8", --30F0
  X"D9", X"E5", X"D9", X"D5", X"EB", X"CD", X"C0", X"30", --30F8
  X"EB", X"38", X"5A", X"E5", X"CD", X"BA", X"2F", X"78", --3100
  X"A7", X"ED", X"62", X"D9", X"E5", X"ED", X"62", X"D9", --3108
  X"06", X"21", X"18", X"11", X"30", X"05", X"19", X"D9", --3110
  X"ED", X"5A", X"D9", X"D9", X"CB", X"1C", X"CB", X"1D", --3118
  X"D9", X"CB", X"1C", X"CB", X"1D", X"D9", X"CB", X"18", --3120
  X"CB", X"19", X"D9", X"CB", X"19", X"1F", X"10", X"E4", --3128
  X"EB", X"D9", X"EB", X"D9", X"C1", X"E1", X"78", X"81", --3130
  X"20", X"01", X"A7", X"3D", X"3F", X"17", X"3F", X"1F", --3138
  X"F2", X"46", X"31", X"30", X"68", X"A7", X"3C", X"20", --3140
  X"08", X"38", X"06", X"D9", X"CB", X"7A", X"D9", X"20", --3148
  X"5C", X"77", X"D9", X"78", X"D9", X"30", X"15", X"7E", --3150
  X"A7", X"3E", X"80", X"28", X"01", X"AF", X"D9", X"A2", --3158
  X"CD", X"FB", X"2F", X"07", X"77", X"38", X"2E", X"23", --3160
  X"77", X"2B", X"18", X"29", X"06", X"20", X"D9", X"CB", --3168
  X"7A", X"D9", X"20", X"12", X"07", X"CB", X"13", X"CB", --3170
  X"12", X"D9", X"CB", X"13", X"CB", X"12", X"D9", X"35", --3178
  X"28", X"D7", X"10", X"EA", X"18", X"D7", X"17", X"30", --3180
  X"0C", X"CD", X"04", X"30", X"20", X"07", X"D9", X"16", --3188
  X"80", X"D9", X"34", X"28", X"18", X"E5", X"23", X"D9", --3190
  X"D5", X"D9", X"C1", X"78", X"17", X"CB", X"16", X"1F", --3198
  X"77", X"23", X"71", X"23", X"72", X"23", X"73", X"E1", --31A0
  X"D1", X"D9", X"E1", X"D9", X"C9", X"CF", X"05", X"CD", --31A8
  X"93", X"32", X"EB", X"AF", X"CD", X"C0", X"30", X"38", --31B0
  X"F4", X"EB", X"CD", X"C0", X"30", X"D8", X"D9", X"E5", --31B8
  X"D9", X"D5", X"E5", X"CD", X"BA", X"2F", X"D9", X"E5", --31C0
  X"60", X"69", X"D9", X"61", X"68", X"AF", X"06", X"DF", --31C8
  X"18", X"10", X"17", X"CB", X"11", X"D9", X"CB", X"11", --31D0
  X"CB", X"10", X"D9", X"29", X"D9", X"ED", X"6A", X"D9", --31D8
  X"38", X"10", X"ED", X"52", X"D9", X"ED", X"52", X"D9", --31E0
  X"30", X"0F", X"19", X"D9", X"ED", X"5A", X"D9", X"A7", --31E8
  X"18", X"08", X"A7", X"ED", X"52", X"D9", X"ED", X"52", --31F0
  X"D9", X"37", X"04", X"FA", X"D2", X"31", X"F5", X"28", --31F8
  X"E1", X"5F", X"51", X"D9", X"59", X"50", X"F1", X"CB", --3200
  X"18", X"F1", X"CB", X"18", X"D9", X"C1", X"E1", X"78", --3208
  X"91", X"C3", X"3D", X"31", X"7E", X"A7", X"C8", X"FE", --3210
  X"81", X"30", X"06", X"36", X"00", X"3E", X"20", X"18", --3218
  X"51", X"FE", X"91", X"20", X"1A", X"23", X"23", X"23", --3220
  X"3E", X"80", X"A6", X"2B", X"B6", X"2B", X"20", X"03", --3228
  X"3E", X"80", X"AE", X"2B", X"20", X"36", X"77", X"23", --3230
  X"36", X"FF", X"2B", X"3E", X"18", X"18", X"33", X"30", --3238
  X"2C", X"D5", X"2F", X"C6", X"91", X"23", X"56", X"23", --3240
  X"5E", X"2B", X"2B", X"0E", X"00", X"CB", X"7A", X"28", --3248
  X"01", X"0D", X"CB", X"FA", X"06", X"08", X"90", X"80", --3250
  X"38", X"04", X"5A", X"16", X"00", X"90", X"28", X"07", --3258
  X"47", X"CB", X"3A", X"CB", X"1B", X"10", X"FA", X"CD", --3260
  X"8E", X"2D", X"D1", X"C9", X"7E", X"D6", X"A0", X"F0", --3268
  X"ED", X"44", X"D5", X"EB", X"2B", X"47", X"CB", X"38", --3270
  X"CB", X"38", X"CB", X"38", X"28", X"05", X"36", X"00", --3278
  X"2B", X"10", X"FB", X"E6", X"07", X"28", X"09", X"47", --3280
  X"3E", X"FF", X"CB", X"27", X"10", X"FC", X"A6", X"77", --3288
  X"EB", X"D1", X"C9", X"CD", X"96", X"32", X"EB", X"7E", --3290
  X"A7", X"C0", X"D5", X"CD", X"7F", X"2D", X"AF", X"23", --3298
  X"77", X"2B", X"77", X"06", X"91", X"7A", X"A7", X"20", --32A0
  X"08", X"B3", X"42", X"28", X"10", X"53", X"58", X"06", --32A8
  X"89", X"EB", X"05", X"29", X"30", X"FC", X"CB", X"09", --32B0
  X"CB", X"1C", X"CB", X"1D", X"EB", X"2B", X"73", X"2B", --32B8
  X"72", X"2B", X"70", X"D1", X"C9", X"00", X"B0", X"00", --32C0
  X"40", X"B0", X"00", X"01", X"30", X"00", X"F1", X"49", --32C8
  X"0F", X"DA", X"A2", X"40", X"B0", X"00", X"0A", X"8F", --32D0
  X"36", X"3C", X"34", X"A1", X"33", X"0F", X"30", X"CA", --32D8
  X"30", X"AF", X"31", X"51", X"38", X"1B", X"35", X"24", --32E0
  X"35", X"3B", X"35", X"3B", X"35", X"3B", X"35", X"3B", --32E8
  X"35", X"3B", X"35", X"3B", X"35", X"14", X"30", X"2D", --32F0
  X"35", X"3B", X"35", X"3B", X"35", X"3B", X"35", X"3B", --32F8
  X"35", X"3B", X"35", X"3B", X"35", X"9C", X"35", X"DE", --3300
  X"35", X"BC", X"34", X"45", X"36", X"6E", X"34", X"69", --3308
  X"36", X"DE", X"35", X"74", X"36", X"B5", X"37", X"AA", --3310
  X"37", X"DA", X"37", X"33", X"38", X"43", X"38", X"E2", --3318
  X"37", X"13", X"37", X"C4", X"36", X"AF", X"36", X"4A", --3320
  X"38", X"92", X"34", X"6A", X"34", X"AC", X"34", X"A5", --3328
  X"34", X"B3", X"34", X"1F", X"36", X"C9", X"35", X"01", --3330
  X"35", X"C0", X"33", X"A0", X"36", X"86", X"36", X"C6", --3338
  X"33", X"7A", X"36", X"06", X"35", X"F9", X"34", X"9B", --3340
  X"36", X"83", X"37", X"14", X"32", X"A2", X"33", X"4F", --3348
  X"2D", X"97", X"32", X"49", X"34", X"1B", X"34", X"2D", --3350
  X"34", X"0F", X"34", X"CD", X"BF", X"35", X"78", X"32", --3358
  X"67", X"5C", X"D9", X"E3", X"D9", X"ED", X"53", X"65", --3360
  X"5C", X"D9", X"7E", X"23", X"E5", X"A7", X"F2", X"80", --3368
  X"33", X"57", X"E6", X"60", X"0F", X"0F", X"0F", X"0F", --3370
  X"C6", X"7C", X"6F", X"7A", X"E6", X"1F", X"18", X"0E", --3378
  X"FE", X"18", X"30", X"08", X"D9", X"01", X"FB", X"FF", --3380
  X"54", X"5D", X"09", X"D9", X"07", X"6F", X"11", X"D7", --3388
  X"32", X"26", X"00", X"19", X"5E", X"23", X"56", X"21", --3390
  X"65", X"33", X"E3", X"D5", X"D9", X"ED", X"4B", X"66", --3398
  X"5C", X"C9", X"F1", X"3A", X"67", X"5C", X"D9", X"18", --33A0
  X"C3", X"D5", X"E5", X"01", X"05", X"00", X"CD", X"05", --33A8
  X"1F", X"E1", X"D1", X"C9", X"ED", X"5B", X"65", X"5C", --33B0
  X"CD", X"C0", X"33", X"ED", X"53", X"65", X"5C", X"C9", --33B8
  X"CD", X"A9", X"33", X"ED", X"B0", X"C9", X"62", X"6B", --33C0
  X"CD", X"A9", X"33", X"D9", X"E5", X"D9", X"E3", X"C5", --33C8
  X"7E", X"E6", X"C0", X"07", X"07", X"4F", X"0C", X"7E", --33D0
  X"E6", X"3F", X"20", X"02", X"23", X"7E", X"C6", X"50", --33D8
  X"12", X"3E", X"05", X"91", X"23", X"13", X"06", X"00", --33E0
  X"ED", X"B0", X"C1", X"E3", X"D9", X"E1", X"D9", X"47", --33E8
  X"AF", X"05", X"C8", X"12", X"13", X"18", X"FA", X"A7", --33F0
  X"C8", X"F5", X"D5", X"11", X"00", X"00", X"CD", X"C8", --33F8
  X"33", X"D1", X"F1", X"3D", X"18", X"F2", X"4F", X"07", --3400
  X"07", X"81", X"4F", X"06", X"00", X"09", X"C9", X"D5", --3408
  X"2A", X"68", X"5C", X"CD", X"06", X"34", X"CD", X"C0", --3410
  X"33", X"E1", X"C9", X"62", X"6B", X"D9", X"E5", X"21", --3418
  X"C5", X"32", X"D9", X"CD", X"F7", X"33", X"CD", X"C8", --3420
  X"33", X"D9", X"E1", X"D9", X"C9", X"E5", X"EB", X"2A", --3428
  X"68", X"5C", X"CD", X"06", X"34", X"EB", X"CD", X"C0", --3430
  X"33", X"EB", X"E1", X"C9", X"06", X"05", X"1A", X"4E", --3438
  X"EB", X"12", X"71", X"23", X"13", X"10", X"F7", X"EB", --3440
  X"C9", X"47", X"CD", X"5E", X"33", X"31", X"0F", X"C0", --3448
  X"02", X"A0", X"C2", X"31", X"E0", X"04", X"E2", X"C1", --3450
  X"03", X"38", X"CD", X"C6", X"33", X"CD", X"62", X"33", --3458
  X"0F", X"01", X"C2", X"02", X"35", X"EE", X"E1", X"03", --3460
  X"38", X"C9", X"06", X"FF", X"18", X"06", X"CD", X"E9", --3468
  X"34", X"D8", X"06", X"00", X"7E", X"A7", X"28", X"0B", --3470
  X"23", X"78", X"E6", X"80", X"B6", X"17", X"3F", X"1F", --3478
  X"77", X"2B", X"C9", X"D5", X"E5", X"CD", X"7F", X"2D", --3480
  X"E1", X"78", X"B1", X"2F", X"4F", X"CD", X"8E", X"2D", --3488
  X"D1", X"C9", X"CD", X"E9", X"34", X"D8", X"D5", X"11", --3490
  X"01", X"00", X"23", X"CB", X"16", X"2B", X"9F", X"4F", --3498
  X"CD", X"8E", X"2D", X"D1", X"C9", X"CD", X"99", X"1E", --34A0
  X"ED", X"78", X"18", X"04", X"CD", X"99", X"1E", X"0A", --34A8
  X"C3", X"28", X"2D", X"CD", X"99", X"1E", X"21", X"2B", --34B0
  X"2D", X"E5", X"C5", X"C9", X"CD", X"F1", X"2B", X"0B", --34B8
  X"78", X"B1", X"20", X"23", X"1A", X"CD", X"8D", X"2C", --34C0
  X"38", X"09", X"D6", X"90", X"38", X"19", X"FE", X"15", --34C8
  X"30", X"15", X"3C", X"3D", X"87", X"87", X"87", X"FE", --34D0
  X"A8", X"30", X"0C", X"ED", X"4B", X"7B", X"5C", X"81", --34D8
  X"4F", X"30", X"01", X"04", X"C3", X"2B", X"2D", X"CF", --34E0
  X"09", X"E5", X"C5", X"47", X"7E", X"23", X"B6", X"23", --34E8
  X"B6", X"23", X"B6", X"78", X"C1", X"E1", X"C0", X"37", --34F0
  X"C9", X"CD", X"E9", X"34", X"D8", X"3E", X"FF", X"18", --34F8
  X"06", X"CD", X"E9", X"34", X"18", X"05", X"AF", X"23", --3500
  X"AE", X"2B", X"07", X"E5", X"3E", X"00", X"77", X"23", --3508
  X"77", X"23", X"17", X"77", X"1F", X"23", X"77", X"23", --3510
  X"77", X"E1", X"C9", X"EB", X"CD", X"E9", X"34", X"EB", --3518
  X"D8", X"37", X"18", X"E7", X"EB", X"CD", X"E9", X"34", --3520
  X"EB", X"D0", X"A7", X"18", X"DE", X"EB", X"CD", X"E9", --3528
  X"34", X"EB", X"D0", X"D5", X"1B", X"AF", X"12", X"1B", --3530
  X"12", X"D1", X"C9", X"78", X"D6", X"08", X"CB", X"57", --3538
  X"20", X"01", X"3D", X"0F", X"30", X"08", X"F5", X"E5", --3540
  X"CD", X"3C", X"34", X"D1", X"EB", X"F1", X"CB", X"57", --3548
  X"20", X"07", X"0F", X"F5", X"CD", X"0F", X"30", X"18", --3550
  X"33", X"0F", X"F5", X"CD", X"F1", X"2B", X"D5", X"C5", --3558
  X"CD", X"F1", X"2B", X"E1", X"7C", X"B5", X"E3", X"78", --3560
  X"20", X"0B", X"B1", X"C1", X"28", X"04", X"F1", X"3F", --3568
  X"18", X"16", X"F1", X"18", X"13", X"B1", X"28", X"0D", --3570
  X"1A", X"96", X"38", X"09", X"20", X"ED", X"0B", X"13", --3578
  X"23", X"E3", X"2B", X"18", X"DF", X"C1", X"F1", X"A7", --3580
  X"F5", X"EF", X"A0", X"38", X"F1", X"F5", X"DC", X"01", --3588
  X"35", X"F1", X"F5", X"D4", X"F9", X"34", X"F1", X"0F", --3590
  X"D4", X"01", X"35", X"C9", X"CD", X"F1", X"2B", X"D5", --3598
  X"C5", X"CD", X"F1", X"2B", X"E1", X"E5", X"D5", X"C5", --35A0
  X"09", X"44", X"4D", X"F7", X"CD", X"B2", X"2A", X"C1", --35A8
  X"E1", X"78", X"B1", X"28", X"02", X"ED", X"B0", X"C1", --35B0
  X"E1", X"78", X"B1", X"28", X"02", X"ED", X"B0", X"2A", --35B8
  X"65", X"5C", X"11", X"FB", X"FF", X"E5", X"19", X"D1", --35C0
  X"C9", X"CD", X"D5", X"2D", X"38", X"0E", X"20", X"0C", --35C8
  X"F5", X"01", X"01", X"00", X"F7", X"F1", X"12", X"CD", --35D0
  X"B2", X"2A", X"EB", X"C9", X"CF", X"0A", X"2A", X"5D", --35D8
  X"5C", X"E5", X"78", X"C6", X"E3", X"9F", X"F5", X"CD", --35E0
  X"F1", X"2B", X"D5", X"03", X"F7", X"E1", X"ED", X"53", --35E8
  X"5D", X"5C", X"D5", X"ED", X"B0", X"EB", X"2B", X"36", --35F0
  X"0D", X"FD", X"CB", X"01", X"BE", X"CD", X"FB", X"24", --35F8
  X"DF", X"FE", X"0D", X"20", X"07", X"E1", X"F1", X"FD", --3600
  X"AE", X"01", X"E6", X"40", X"C2", X"8A", X"1C", X"22", --3608
  X"5D", X"5C", X"FD", X"CB", X"01", X"FE", X"CD", X"FB", --3610
  X"24", X"E1", X"22", X"5D", X"5C", X"18", X"A0", X"01", --3618
  X"01", X"00", X"F7", X"22", X"5B", X"5C", X"E5", X"2A", --3620
  X"51", X"5C", X"E5", X"3E", X"FF", X"CD", X"01", X"16", --3628
  X"CD", X"E3", X"2D", X"E1", X"CD", X"15", X"16", X"D1", --3630
  X"2A", X"5B", X"5C", X"A7", X"ED", X"52", X"44", X"4D", --3638
  X"CD", X"B2", X"2A", X"EB", X"C9", X"CD", X"94", X"1E", --3640
  X"FE", X"10", X"D2", X"9F", X"1E", X"2A", X"51", X"5C", --3648
  X"E5", X"CD", X"01", X"16", X"CD", X"E6", X"15", X"01", --3650
  X"00", X"00", X"30", X"03", X"0C", X"F7", X"12", X"CD", --3658
  X"B2", X"2A", X"E1", X"CD", X"15", X"16", X"C3", X"BF", --3660
  X"35", X"CD", X"F1", X"2B", X"78", X"B1", X"28", X"01", --3668
  X"1A", X"C3", X"28", X"2D", X"CD", X"F1", X"2B", X"C3", --3670
  X"2B", X"2D", X"D9", X"E5", X"21", X"67", X"5C", X"35", --3678
  X"E1", X"20", X"04", X"23", X"D9", X"C9", X"D9", X"5E", --3680
  X"7B", X"17", X"9F", X"57", X"19", X"D9", X"C9", X"13", --3688
  X"13", X"1A", X"1B", X"1B", X"A7", X"20", X"EF", X"D9", --3690
  X"23", X"D9", X"C9", X"F1", X"D9", X"E3", X"D9", X"C9", --3698
  X"EF", X"C0", X"02", X"31", X"E0", X"05", X"27", X"E0", --36A0
  X"01", X"C0", X"04", X"03", X"E0", X"38", X"C9", X"EF", --36A8
  X"31", X"36", X"00", X"04", X"3A", X"38", X"C9", X"31", --36B0
  X"3A", X"C0", X"03", X"E0", X"01", X"30", X"00", X"03", --36B8
  X"A1", X"03", X"38", X"C9", X"EF", X"3D", X"34", X"F1", --36C0
  X"38", X"AA", X"3B", X"29", X"04", X"31", X"27", X"C3", --36C8
  X"03", X"31", X"0F", X"A1", X"03", X"88", X"13", X"36", --36D0
  X"58", X"65", X"66", X"9D", X"78", X"65", X"40", X"A2", --36D8
  X"60", X"32", X"C9", X"E7", X"21", X"F7", X"AF", X"24", --36E0
  X"EB", X"2F", X"B0", X"B0", X"14", X"EE", X"7E", X"BB", --36E8
  X"94", X"58", X"F1", X"3A", X"7E", X"F8", X"CF", X"E3", --36F0
  X"38", X"CD", X"D5", X"2D", X"20", X"07", X"38", X"03", --36F8
  X"86", X"30", X"09", X"CF", X"05", X"38", X"07", X"96", --3700
  X"30", X"04", X"ED", X"44", X"77", X"C9", X"EF", X"02", --3708
  X"A0", X"38", X"C9", X"EF", X"3D", X"31", X"37", X"00", --3710
  X"04", X"38", X"CF", X"09", X"A0", X"02", X"38", X"7E", --3718
  X"36", X"80", X"CD", X"28", X"2D", X"EF", X"34", X"38", --3720
  X"00", X"03", X"01", X"31", X"34", X"F0", X"4C", X"CC", --3728
  X"CC", X"CD", X"03", X"37", X"00", X"08", X"01", X"A1", --3730
  X"03", X"01", X"38", X"34", X"EF", X"01", X"34", X"F0", --3738
  X"31", X"72", X"17", X"F8", X"04", X"01", X"A2", X"03", --3740
  X"A2", X"03", X"31", X"34", X"32", X"20", X"04", X"A2", --3748
  X"03", X"8C", X"11", X"AC", X"14", X"09", X"56", X"DA", --3750
  X"A5", X"59", X"30", X"C5", X"5C", X"90", X"AA", X"9E", --3758
  X"70", X"6F", X"61", X"A1", X"CB", X"DA", X"96", X"A4", --3760
  X"31", X"9F", X"B4", X"E7", X"A0", X"FE", X"5C", X"FC", --3768
  X"EA", X"1B", X"43", X"CA", X"36", X"ED", X"A7", X"9C", --3770
  X"7E", X"5E", X"F0", X"6E", X"23", X"80", X"93", X"04", --3778
  X"0F", X"38", X"C9", X"EF", X"3D", X"34", X"EE", X"22", --3780
  X"F9", X"83", X"6E", X"04", X"31", X"A2", X"0F", X"27", --3788
  X"03", X"31", X"0F", X"31", X"0F", X"31", X"2A", X"A1", --3790
  X"03", X"31", X"37", X"C0", X"00", X"04", X"02", X"38", --3798
  X"C9", X"A1", X"03", X"01", X"36", X"00", X"02", X"1B", --37A0
  X"38", X"C9", X"EF", X"39", X"2A", X"A1", X"03", X"E0", --37A8
  X"00", X"06", X"1B", X"33", X"03", X"EF", X"39", X"31", --37B0
  X"31", X"04", X"31", X"0F", X"A1", X"03", X"86", X"14", --37B8
  X"E6", X"5C", X"1F", X"0B", X"A3", X"8F", X"38", X"EE", --37C0
  X"E9", X"15", X"63", X"BB", X"23", X"EE", X"92", X"0D", --37C8
  X"CD", X"ED", X"F1", X"23", X"5D", X"1B", X"EA", X"04", --37D0
  X"38", X"C9", X"EF", X"31", X"1F", X"01", X"20", X"05", --37D8
  X"38", X"C9", X"CD", X"97", X"32", X"7E", X"FE", X"81", --37E0
  X"38", X"0E", X"EF", X"A1", X"1B", X"01", X"05", X"31", --37E8
  X"36", X"A3", X"01", X"00", X"06", X"1B", X"33", X"03", --37F0
  X"EF", X"A0", X"01", X"31", X"31", X"04", X"31", X"0F", --37F8
  X"A1", X"03", X"8C", X"10", X"B2", X"13", X"0E", X"55", --3800
  X"E4", X"8D", X"58", X"39", X"BC", X"5B", X"98", X"FD", --3808
  X"9E", X"00", X"36", X"75", X"A0", X"DB", X"E8", X"B4", --3810
  X"63", X"42", X"C4", X"E6", X"B5", X"09", X"36", X"BE", --3818
  X"E9", X"36", X"73", X"1B", X"5D", X"EC", X"D8", X"DE", --3820
  X"63", X"BE", X"F0", X"61", X"A1", X"B3", X"0C", X"04", --3828
  X"0F", X"38", X"C9", X"EF", X"31", X"31", X"04", X"A1", --3830
  X"03", X"1B", X"28", X"A1", X"0F", X"05", X"24", X"31", --3838
  X"0F", X"38", X"C9", X"EF", X"22", X"A3", X"03", X"1B", --3840
  X"38", X"C9", X"EF", X"31", X"30", X"00", X"1E", X"A2", --3848
  X"38", X"EF", X"01", X"31", X"30", X"00", X"07", X"25", --3850
  X"04", X"38", X"C3", X"C4", X"36", X"02", X"31", X"30", --3858
  X"00", X"09", X"A0", X"01", X"37", X"00", X"06", X"A1", --3860
  X"01", X"05", X"02", X"A1", X"38", X"C9", X"FF", X"FF", --3868
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3870
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3878
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3880
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3888
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3890
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3898
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --38F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3900
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3908
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3910
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3918
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3920
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3928
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3930
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3938
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3940
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3948
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3950
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3958
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3960
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3968
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3970
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3978
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3980
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3988
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3990
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3998
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39A0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39A8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39B0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39B8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39C0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39C8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39D0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39D8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39E0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39E8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39F0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --39F8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3A98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3AF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3B98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3BF8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C00
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C08
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C10
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C18
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C20
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C28
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C30
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C38
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C40
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C48
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C50
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C58
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C60
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C68
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C70
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C78
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C80
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C88
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C90
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3C98
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CA0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CA8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CB0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CB8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CC0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CC8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CD0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CD8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CE0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CE8
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CF0
  X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", --3CF8
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", --3D00
  X"00", X"10", X"10", X"10", X"10", X"00", X"10", X"00", --3D08
  X"00", X"24", X"24", X"00", X"00", X"00", X"00", X"00", --3D10
  X"00", X"24", X"7E", X"24", X"24", X"7E", X"24", X"00", --3D18
  X"00", X"08", X"3E", X"28", X"3E", X"0A", X"3E", X"08", --3D20
  X"00", X"62", X"64", X"08", X"10", X"26", X"46", X"00", --3D28
  X"00", X"10", X"28", X"10", X"2A", X"44", X"3A", X"00", --3D30
  X"00", X"08", X"10", X"00", X"00", X"00", X"00", X"00", --3D38
  X"00", X"04", X"08", X"08", X"08", X"08", X"04", X"00", --3D40
  X"00", X"20", X"10", X"10", X"10", X"10", X"20", X"00", --3D48
  X"00", X"00", X"14", X"08", X"3E", X"08", X"14", X"00", --3D50
  X"00", X"00", X"08", X"08", X"3E", X"08", X"08", X"00", --3D58
  X"00", X"00", X"00", X"00", X"00", X"08", X"08", X"10", --3D60
  X"00", X"00", X"00", X"00", X"3E", X"00", X"00", X"00", --3D68
  X"00", X"00", X"00", X"00", X"00", X"18", X"18", X"00", --3D70
  X"00", X"00", X"02", X"04", X"08", X"10", X"20", X"00", --3D78
  X"00", X"3C", X"46", X"4A", X"52", X"62", X"3C", X"00", --3D80
  X"00", X"18", X"28", X"08", X"08", X"08", X"3E", X"00", --3D88
  X"00", X"3C", X"42", X"02", X"3C", X"40", X"7E", X"00", --3D90
  X"00", X"3C", X"42", X"0C", X"02", X"42", X"3C", X"00", --3D98
  X"00", X"08", X"18", X"28", X"48", X"7E", X"08", X"00", --3DA0
  X"00", X"7E", X"40", X"7C", X"02", X"42", X"3C", X"00", --3DA8
  X"00", X"3C", X"40", X"7C", X"42", X"42", X"3C", X"00", --3DB0
  X"00", X"7E", X"02", X"04", X"08", X"10", X"10", X"00", --3DB8
  X"00", X"3C", X"42", X"3C", X"42", X"42", X"3C", X"00", --3DC0
  X"00", X"3C", X"42", X"42", X"3E", X"02", X"3C", X"00", --3DC8
  X"00", X"00", X"00", X"10", X"00", X"00", X"10", X"00", --3DD0
  X"00", X"00", X"10", X"00", X"00", X"10", X"10", X"20", --3DD8
  X"00", X"00", X"04", X"08", X"10", X"08", X"04", X"00", --3DE0
  X"00", X"00", X"00", X"3E", X"00", X"3E", X"00", X"00", --3DE8
  X"00", X"00", X"10", X"08", X"04", X"08", X"10", X"00", --3DF0
  X"00", X"3C", X"42", X"04", X"08", X"00", X"08", X"00", --3DF8
  X"00", X"3C", X"4A", X"56", X"5E", X"40", X"3C", X"00", --3E00
  X"00", X"3C", X"42", X"42", X"7E", X"42", X"42", X"00", --3E08
  X"00", X"7C", X"42", X"7C", X"42", X"42", X"7C", X"00", --3E10
  X"00", X"3C", X"42", X"40", X"40", X"42", X"3C", X"00", --3E18
  X"00", X"78", X"44", X"42", X"42", X"44", X"78", X"00", --3E20
  X"00", X"7E", X"40", X"7C", X"40", X"40", X"7E", X"00", --3E28
  X"00", X"7E", X"40", X"7C", X"40", X"40", X"40", X"00", --3E30
  X"00", X"3C", X"42", X"40", X"4E", X"42", X"3C", X"00", --3E38
  X"00", X"42", X"42", X"7E", X"42", X"42", X"42", X"00", --3E40
  X"00", X"3E", X"08", X"08", X"08", X"08", X"3E", X"00", --3E48
  X"00", X"02", X"02", X"02", X"42", X"42", X"3C", X"00", --3E50
  X"00", X"44", X"48", X"70", X"48", X"44", X"42", X"00", --3E58
  X"00", X"40", X"40", X"40", X"40", X"40", X"7E", X"00", --3E60
  X"00", X"42", X"66", X"5A", X"42", X"42", X"42", X"00", --3E68
  X"00", X"42", X"62", X"52", X"4A", X"46", X"42", X"00", --3E70
  X"00", X"3C", X"42", X"42", X"42", X"42", X"3C", X"00", --3E78
  X"00", X"7C", X"42", X"42", X"7C", X"40", X"40", X"00", --3E80
  X"00", X"3C", X"42", X"42", X"52", X"4A", X"3C", X"00", --3E88
  X"00", X"7C", X"42", X"42", X"7C", X"44", X"42", X"00", --3E90
  X"00", X"3C", X"40", X"3C", X"02", X"42", X"3C", X"00", --3E98
  X"00", X"FE", X"10", X"10", X"10", X"10", X"10", X"00", --3EA0
  X"00", X"42", X"42", X"42", X"42", X"42", X"3C", X"00", --3EA8
  X"00", X"42", X"42", X"42", X"42", X"24", X"18", X"00", --3EB0
  X"00", X"42", X"42", X"42", X"42", X"5A", X"24", X"00", --3EB8
  X"00", X"42", X"24", X"18", X"18", X"24", X"42", X"00", --3EC0
  X"00", X"82", X"44", X"28", X"10", X"10", X"10", X"00", --3EC8
  X"00", X"7E", X"04", X"08", X"10", X"20", X"7E", X"00", --3ED0
  X"00", X"0E", X"08", X"08", X"08", X"08", X"0E", X"00", --3ED8
  X"00", X"00", X"40", X"20", X"10", X"08", X"04", X"00", --3EE0
  X"00", X"70", X"10", X"10", X"10", X"10", X"70", X"00", --3EE8
  X"00", X"10", X"38", X"54", X"10", X"10", X"10", X"00", --3EF0
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"FF", --3EF8
  X"00", X"1C", X"22", X"78", X"20", X"20", X"7E", X"00", --3F00
  X"00", X"00", X"38", X"04", X"3C", X"44", X"3C", X"00", --3F08
  X"00", X"20", X"20", X"3C", X"22", X"22", X"3C", X"00", --3F10
  X"00", X"00", X"1C", X"20", X"20", X"20", X"1C", X"00", --3F18
  X"00", X"04", X"04", X"3C", X"44", X"44", X"3C", X"00", --3F20
  X"00", X"00", X"38", X"44", X"78", X"40", X"3C", X"00", --3F28
  X"00", X"0C", X"10", X"18", X"10", X"10", X"10", X"00", --3F30
  X"00", X"00", X"3C", X"44", X"44", X"3C", X"04", X"38", --3F38
  X"00", X"40", X"40", X"78", X"44", X"44", X"44", X"00", --3F40
  X"00", X"10", X"00", X"30", X"10", X"10", X"38", X"00", --3F48
  X"00", X"04", X"00", X"04", X"04", X"04", X"24", X"18", --3F50
  X"00", X"20", X"28", X"30", X"30", X"28", X"24", X"00", --3F58
  X"00", X"10", X"10", X"10", X"10", X"10", X"0C", X"00", --3F60
  X"00", X"00", X"68", X"54", X"54", X"54", X"54", X"00", --3F68
  X"00", X"00", X"78", X"44", X"44", X"44", X"44", X"00", --3F70
  X"00", X"00", X"38", X"44", X"44", X"44", X"38", X"00", --3F78
  X"00", X"00", X"78", X"44", X"44", X"78", X"40", X"40", --3F80
  X"00", X"00", X"3C", X"44", X"44", X"3C", X"04", X"06", --3F88
  X"00", X"00", X"1C", X"20", X"20", X"20", X"20", X"00", --3F90
  X"00", X"00", X"38", X"40", X"38", X"04", X"78", X"00", --3F98
  X"00", X"10", X"38", X"10", X"10", X"10", X"0C", X"00", --3FA0
  X"00", X"00", X"44", X"44", X"44", X"44", X"38", X"00", --3FA8
  X"00", X"00", X"44", X"44", X"28", X"28", X"10", X"00", --3FB0
  X"00", X"00", X"44", X"54", X"54", X"54", X"28", X"00", --3FB8
  X"00", X"00", X"44", X"28", X"10", X"28", X"44", X"00", --3FC0
  X"00", X"00", X"44", X"44", X"44", X"3C", X"04", X"38", --3FC8
  X"00", X"00", X"7C", X"08", X"10", X"20", X"7C", X"00", --3FD0
  X"00", X"0E", X"08", X"30", X"08", X"08", X"0E", X"00", --3FD8
  X"00", X"08", X"08", X"08", X"08", X"08", X"08", X"00", --3FE0
  X"00", X"70", X"10", X"0C", X"10", X"10", X"70", X"00", --3FE8
  X"00", X"14", X"28", X"00", X"00", X"00", X"00", X"00", --3FF0
  X"3C", X"42", X"99", X"A1", X"A1", X"99", X"42", X"3C");--3FF8

begin

  process (clk)
  begin
    if rising_edge(clk) then
      dout <= rom(to_integer(unsigned(addr)));
    end if;
  end process;

end behavioral;
