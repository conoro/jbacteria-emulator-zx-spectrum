library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

entity vram is port(
    clk     : in  std_logic;
    addr    : in  std_logic_vector(13 downto 0);
    dataout : out std_logic_vector( 7 downto 0));
end vram;

architecture Behavioral of vram is

  type arrayen is array(3 downto 0) of std_logic;
  type arraydo is array(3 downto 0) of std_logic_vector(7 downto 0);
  signal en : arrayen;
  signal do : arraydo;

begin
  process(addr, do)
  variable i : integer;
  begin
    dataout <= (others => '0');
    for i in 0 to 3 loop
      en(i) <= '0';
      if (to_integer(unsigned(addr(13 downto 11))) = i) then
        en(i) <= '1';
        dataout <= do(i);
      end if;
    end loop;
  end process;

  ram0 : RAMB16_S9
  generic map (
      write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    , INIT_00   => X"579500912A0140F5FFFFFFFF7CF003E00FE50BE080B8FFBFAAAA9057550A0000"
    , INIT_01   => X"FF5F155F55FF55555555FFFFDC035EF5100206F8A1E1F72B480000FFFF561000"
    , INIT_02   => X"5D005715D5D4D45F55FF7F7F136FFD7F0C6DFCFF80E2FC0B00AAFFB4F7572100"
    , INIT_03   => X"5500AA8201D5FFFFFF0B0010D4870055850AFD00DF10F4400A8055F5FB570900"
    , INIT_04   => X"5F5505411540EA004080000815F957AF5C1502F40711D100AFFDFFFF5E250000"
    , INIT_05   => X"551555D5FF5F40150055EF7DD1FD571DFB3F94F5061C77AB5751552102020000"
    , INIT_06   => X"550000D4DDFE3FD5BF852254A1F3FF97F8757FDEE24100005F55440001000000"
    , INIT_07   => X"5509020800D5FF630E3CC2FFBF11585EDFDFFE9F300997F0D595142400000000"
    , INIT_08   => X"BF2A0044550080AAF7FFFF7F3EFC07B407DA1DF0200CFF5D415505FDAA800000"
    , INIT_09   => X"BFAA02FFABEBAAEFAE2AFF7F6C8FFFCF2981EBFF5FE1E70715804AEFFF0B0500"
    , INIT_0A   => X"2B00AA0AAA68F8FFAFFF5F1F099E7C002C2E00FC00F1FE150050FDEAFE3D0000"
    , INIT_0B   => X"2A015429AAFAFFFF7F040088EACB00BE0220EA80DF08EC105520AA7FFF2F0000"
    , INIT_0C   => X"FFAA28A8AAA85C0A004280885AFC8B5EAFEA2920E623B32055EEFFAFAB8A0000"
    , INIT_0D   => X"AFA2A0AADAFB00B004ABEEFF90FBAB2DFEFF29F10438FF45AF8AAA8A08000000"
    , INIT_0E   => X"AA0000A8AAEB7FF87FAD148000B95E2D78EF1EBFA3838200B702000000000000"
    , INIT_0F   => X"AA000000147AFF4F3E04E257FF10B3B87FDDFD1D28118BB0AA2A400000000000"
    , INIT_10   => X"FF5705902A0009F5FE7FED3F1B8E0DF413B51FF8C831FE2F800A20BF57250000"
    , INIT_11   => X"FF57155755FD55555555FF1F2CFCFFFF13C2FDFFBFC1E70A2A2900FDFF560000"
    , INIT_12   => X"9540551545D0B47F55FF2F1F04FD00000DAD00808072FC4B00A8FFB4FB5F0900"
    , INIT_13   => X"5704A10255F5FFFF23060044F5C5007D0540D940DF10E8402A007FEBFF550400"
    , INIT_14   => X"5F55455155D5F0818056545059FC17F95100D6C0F012B580AF55757555200000"
    , INIT_15   => X"551500D57FFF4055215FEF7F38FB551DFCFF6D7304707F8B5F55512180000000"
    , INIT_16   => X"1500005455FFFFF1FFF53D408051F5577CED8239874205085E55110200000000"
    , INIT_17   => X"55A508002AD4FF7F6A08F9EBFF99D471FFCF3B9E171395F05155118804000000"
    , INIT_18   => X"BFAA00049500A0AAFFED7FBF1B8739F413FA1FAE86B2FC5600A000FFAD800000"
    , INIT_19   => X"D7AA00BFAAEAFAFFAB22FF0F5CF8B7FF2341BFFD77C1E7075D4055FFFF0B1100"
    , INIT_1A   => X"2A000A0A82E8EAFF2FFF030F02FE01002FEE08000FF9FF1700507FEAFE370000"
    , INIT_1B   => X"2A010400ABFA1F02100200ACFEC303BA0800A080CF08E8005740DABFFFAB0000"
    , INIT_1C   => X"FFABAAAAFFEACC2EA4D6AAB89AFE2B710000AC6BF127B31055BAAFAB2A050000"
    , INIT_1D   => X"AB0840A8F6F701B00AFF97BF7CFE8A2E0400E66B0828FF07BF00040411000000"
    , INIT_1E   => X"AA0000A8AAFA7FE3BFF57120F891AA2ADC6D827DC1848B10AB0A040000000000"
    , INIT_1F   => X"AA0AA0005CEAFFFFD609FFFFFF8809EBDE6B0AB60F128BB0A40A040140000000"
    , INIT_20   => X"EF5F155000005455B5BFD59F97E3F13F34FDFDD71094F92B000400FF5F150200"
    , INIT_21   => X"7F55055555B554555505FF07B8E1E7FB13621F9FB7C1F302BEAAAA6BFF560400"
    , INIT_22   => X"15A0051445B0FCFF55FF2107413D41010FED54007F7CFC2B01A0FAB4FF5F0500"
    , INIT_23   => X"5F049080D7FF07001002C055FFE50F54104050C4EF10D900AA00FFFDFF150000"
    , INIT_24   => X"5F5D55F5AA75305081905D5533FF57E20000589DF917F544AA55555505100000"
    , INIT_25   => X"551500F5BFFF4365558F905F7F5DC51FF8FFE3EF09507F835F55514100000000"
    , INIT_26   => X"5500001545EF7FCD3F1B3D90FF11545F7C6F81F7410405A8D555410000000000"
    , INIT_27   => X"555455053E74FF7F0A1EFFFFFF480AF6DD2F0AF7072247F05151412000000000"
    , INIT_28   => X"BFAA02002A00A9EAFEEAAA9E971B029F05FAF08A2AD8FB17000000FFF7420000"
    , INIT_29   => X"AB2A00AB00EAF8FFAB00FF037042FFFF2721FEFFD3C3F3175D4055FEFF2F1000"
    , INIT_2A   => X"4A000A2A8AE8FAFFAFFF0083A01EAA0A2DEEA800FF7EF85708485FEAFBAF0000"
    , INIT_2B   => X"AB1000007FFD0301100238E9F7E23FA82A00A0A8EF08D90057006DFFFF2A0500"
    , INIT_2C   => X"FFABAAAAFF7E00A72AA7BEBA57FF2FC6F92F30FA7B2FBBA855AAAAAAAA020000"
    , INIT_2D   => X"2A0200A8EAFF07A8AAB3CFFFAFAA384F0800F0EF09A0FF17BF00000812000000"
    , INIT_2E   => X"2A8A0028A0FAFF3C1F6B0EF8D711A836DE4DA1B7A1068B50EA2B101200000000"
    , INIT_2F   => X"AA228A025CEAFFFFFEB3FEDFFFC8047C3B268EF3002668F0040410080A000000"
    , INIT_30   => X"FF5F1500000054555555159DFF01023001FD58C017E9F32B000000FF7F150100"
    , INIT_31   => X"7F85001500D4D45B5505FF01C08DFF7F1622FCFFFFEDF903AAAAFEB5FF5B0100"
    , INIT_32   => X"1740055455D4ECFF5F3F2041501F741505AC5000DF6FF4AF02A0FAF5FE5B1500"
    , INIT_33   => X"5F050000FFFF0300700206F96DF17F00558102D4E710D180BB00FFFFFF150000"
    , INIT_34   => X"555555FDFA5B007755A5E5D5A5FE5786FFFF7BED7B1FF7D2A855555501000000"
    , INIT_35   => X"57010054BFFE0F65D5BCC7FF0755071BE898FDDF7140FFAB6F55840000000000"
    , INIT_36   => X"5500408242F5FF7A0E7A04BEAAF151637E5FD3BF600E97A8F557050000000000"
    , INIT_37   => X"5555511528B4FFFFFE3FFFF7FF4863583B164AF90024317050A1848240000000"
    , INIT_38   => X"FFAA02001400AAAABBAA029AFF01046008FA0C402BF1F305000000FFDF0B0400"
    , INIT_39   => X"AA12000A006A78FFAB00FF00A69301202711010000F1FC2614505DEAFE2F0400"
    , INIT_3A   => X"2B000AAAEFEAFEFFFF1F0020A88FA8AA0848A000FF77F45F555055DAFF2F0000"
    , INIT_3B   => X"ABAA0000FFFF0100400001FEF5F0FFA0AA4205E81728D3005500FFFFFF8A0200"
    , INIT_3C   => X"FFAAAAEAFF7F00F7AF3AFFFACAFDAF0E0380FFEE832EBBFC50AAAA8A48000000"
    , INIT_3D   => X"AA0A00A0EAFB1FE87F9662BA03C8012E5867FEDFF2A1FFD7BF02112200000000"
    , INIT_3E   => X"AA00000090FAFF75004602FFFF11AEBAFF5DFF9F700A8B50EA2B800000000000"
    , INIT_3F   => X"AA8AAA0800EAFFFFFE3FF5E39F48B2507716F4FF00E41EF00404202010080000"
  )
  port map (
      DI    => "00000000"
    , DIP   => "0"
    , DO    => do(0)
    , ADDR  => addr(10 downto 0)
    , CLK   => clk
    , EN    => en(0)
    , WE    => '0'
    , SSR   => '0'
  );

  ram1 : RAMB16_S9
  generic map (
      write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    , INIT_00   => X"5555545540B5FFFFEE3FFAA33F885153EFA8000000CC21F0A150858A04010000"
    , INIT_01   => X"F77F5555BFFFFFFF1B00E0AFFAFFC1C0FFED2EF037C20FFF0000500000950800"
    , INIT_02   => X"FFFFFDFFFFFFFFFFFFC1FF05A8FFF0F9B601F89014E0ED03F8FF0F803F000A00"
    , INIT_03   => X"FFFFFF5F07800700FCE0FF7DE800C4FD56FE632F1720030F06CFFD0FA2AA4300"
    , INIT_04   => X"FFFF1F0055557C0056ED0380801640EED50CF8E00100C13795C07F00AAF63900"
    , INIT_05   => X"FFC038465184FF1F44D5EBA7FFFFE0FCDFACF740005940FF5F0900AA2AAA2001"
    , INIT_06   => X"B7DF5FFDF9BFA87FFF10FDF3037CFEFD47FF2FBB0B017444000A5000B88A4201"
    , INIT_07   => X"0A00D72850C1AF1F7C3FF02AD5FFAFAC0780BB40217047910300000000000000"
    , INIT_08   => X"AAAAAA22AAFAFFFFFC3F52FF0388E136EF08802080C813F80002102050000000"
    , INIT_09   => X"5DABAEEAEAFFFFFF07A07F55D5FFF3EEFF6A976829C40FFE0000EA00002A0000"
    , INIT_0A   => X"FFFFEFFFFFFFC1FFEA81AB02D0FFE8E9AD01FCA024E4CB03E2FFFF01F4032100"
    , INIT_0B   => X"FFFFFF5F0F000700EE403FAFF4008AE94C0605370A40820F0BCFEA070D550200"
    , INIT_0C   => X"FFFF0140A0AA7A00A6FE074050AB00EC5B147FC93000E0370A843E1455BD5C00"
    , INIT_0D   => X"FFE870CC02E1D70F10BADB0FD5FFFCCEFF1CEF4400E480AAAB02005C55445100"
    , INIT_0E   => X"7FF7BFDE5FD5D07FFF109383FF03FFEF011C18411700F0200005000050450100"
    , INIT_0F   => X"1504AF10A4F0D70FF81D78F7EAFF95EC0B40FF0714A107A30300000000000000"
    , INIT_10   => X"5555555551D5FFFFED3F347E0008C1B9DF0855E0408803F88890445505440000"
    , INIT_11   => X"F7FF7557BFFFFFFFE7FFDE026AFFFFF3EFCDC2180CC41FFE0000D40000970200"
    , INIT_12   => X"FFFFFFFFFF0F000FD0030000A8FFF0F9B601FCA024C0CB060DFEFF1FA03F0B00"
    , INIT_13   => X"FFFFFF2F10000F00D640D357EA00C5ECD5AA8E3F2F20821F01CFD4037A000000"
    , INIT_14   => X"FFFF1F005555FC0056D507A8EA5540EED50CBFC4D983E82F55011C00AAEA2E00"
    , INIT_15   => X"FFF5E1980BF8A00F40D5EB0F00FCE7CCEBAC7F0110F800BD5F9500B8AAA02800"
    , INIT_16   => X"EB5F7FFDFFAEE8FFFF10010F00E0EF6D00030E0068A0F06401020008A0A25001"
    , INIT_17   => X"2A105F3011FCEF07B017B8FAFFAF82FC0590774FA0810FC20300000000000000"
    , INIT_18   => X"AEAAAAAAAAFEFFFF7D1D280CE03F81E7BF08AA703F8903FC000010A82A110000"
    , INIT_19   => X"FF76AFBAEAFFFFFF6F75AC01D4FF3FE1FFD0E1E80BC41F1E0000E900002B2000"
    , INIT_1A   => X"FFFFFFFF7F005000A0070000D0FFF8E9AD03FE2245D08F869AF0FF7F447D0200"
    , INIT_1B   => X"FFFFFFCF07F00F00A680AEABF48082E948569DEF5A80801F22CFA802FDC33F00"
    , INIT_1C   => X"FF1F7C00A8AAFA01A3FE4F7DB50A00EE7FFC9FD2E807E46F2B00195554351F04"
    , INIT_1D   => X"7FFAC13D03FED01F10B8FB1FC01FF88EFF5C7F0030F081AAB782007055511400"
    , INIT_1E   => X"57FFBF5A5555F4FFFE90007E00FED5AFC0018500C084E1280101000040450400"
    , INIT_1F   => X"0544AF6101FFDF07E81A58F5FF5580F802C03FE781050FC2010000C0FF3F1E00"
    , INIT_20   => X"D55F555555F5FFFF7D1F4803FF7FC11FBF08FFF01F8B07FE0052425555440000"
    , INIT_21   => X"DFDFFA57DFFEFFFFDF2A5401A8FF3FFDD6D0E24809E01E0E0E00F40000570500"
    , INIT_22   => X"FFFFFFFF03000000C0072000E8FFD0F95603FE5030A08F068DC7FF3F10AA2100"
    , INIT_23   => X"FFFFFFEF1FFF1F00D680FE1FFA40C1ECD50AF88F0040813F08CF5401EAEFFF01"
    , INIT_24   => X"FFFFF1185555FC8149D59F825F5540ECD5FC8FD2C00FEA6F55050380A82A0B01"
    , INIT_25   => X"FFFDC37B80FFA01F40D5D9F37F809FECFBACBF1808F000A55FC500E0AA2A2A00"
    , INIT_26   => X"AB7F7DF4BFABFAFF0ED3008CFFFFEAAD7000A600001EE0500101000080225100"
    , INIT_27   => X"2B105FC283FFBF03701728A8BF2A805C01A04FF7071A1CC6A1010080FF7F3C00"
    , INIT_28   => X"BBAAAAAAEAFFFFFF793E90F0FFFF82FDF8083FB41F8A07FF000028AAAA100000"
    , INIT_29   => X"FFFF5FFDF5FFFFFF7F01A803D0FE1FF9FB70F15012C81E07FD00AA0000BF1000"
    , INIT_2A   => X"FFFFFF7F01000100900FF800D0FFA8E96503FED90F90878646CDFF1F80400701"
    , INIT_2B   => X"FFFFFFFFFFBF3E00A600FC0BF5A080ED58FCCFEF0240C11F02CF2800F5FF1F00"
    , INIT_2C   => X"FF57C7A9AAAAFAC3A0BA7FF8AF0240EEFF14C7DBA00FB46E2B00075541950504"
    , INIT_2D   => X"7FFA8F75C0FFD03F10B8F94301F003FEFFDE1F7C50E0064AFFEA008057151400"
    , INIT_2E   => X"57FFFB785555FDFF007FC004A07FF5AD3800F388006E64A80300000000110400"
    , INIT_2F   => X"0740BE05C2FFFE03E82A0850570580AE00C853C3173808C60106000000000000"
    , INIT_30   => X"EF7F5555BDFEFFFFFB1E201EF8FFC38A471800FA0FC607FF008040F557450200"
    , INIT_31   => X"FFFFF657BFFFFFFFFF20FC07A8FF2FF9D691F15012E81D0FFA0FD53000574500"
    , INIT_32   => X"FFFFFFBF00800300C00FFF5FE8FFD4E9567FFED850A8070F028AFF1F00A41300"
    , INIT_33   => X"FFFFFF5F7D553D0056005185FA5041ECD504F0EF0580C23729CF1000AAFFEF00"
    , INIT_34   => X"FFAB8E335555FC6344D5FBFF551440CCDDFCE7DF402FC07F5F15138282CA0201"
    , INIT_35   => X"BFFF57FFE0FFA03F8052D947813FF0BEFEBEDFF7E0401B445FF54000AE2A0A04"
    , INIT_36   => X"2AFFF5B1AA80FE7F007FE00350BFFEAD1D80FA1403F648D00300000000081100"
    , INIT_37   => X"13107D0AE3FFFD01501518802A00805701A0D1013B00208E010C00F0FF1F0700"
    , INIT_38   => X"BEAAABAAEAFFFFFFFB2FA003D5FFE7C5FF1800F907820FFF0020A4DABE0A0000"
    , INIT_39   => X"FFFFBFFEFBFFFFFFFFA0FE03D0FF1FE9EDE1F89012E87D70F5FFFBFC01AF0000"
    , INIT_3A   => X"FFFFFF5F06800300F01FF7FFD4FFA8E964FF7DD82F50070F00C4FF0F00000700"
    , INIT_3B   => X"FFFFFF81AAAA7E00A6002B00FDAC80EC59FCFFEF0280C037029F0000D5FD7300"
    , INIT_3C   => X"FF5F1CC7A82AFE3790BAFFFFAA0240FEFFFCF7DF8036A0FAAB02095515654100"
    , INIT_3D   => X"7FF5AFD6F1D7D07F0090F9FF7F8078D5FCFE6F7BC1002D4AFFFA20005C150500"
    , INIT_3E   => X"17F7EB6B058AFF3F013F7005A8FFFFAC0F007BAA0CF042A10300000000440400"
    , INIT_3F   => X"0540FA15F7FFFF01A82A1800050080AB00D0A900D83E008F011000E0FF3F0E00"
  )
  port map (
      DI    => "00000000"
    , DIP   => "0"
    , DO    => do(1)
    , ADDR  => addr(10 downto 0)
    , CLK   => clk
    , EN    => en(1)
    , WE    => '0'
    , SSR   => '0'
  );

  ram2 : RAMB16_S9
  generic map (
      write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    , INIT_00   => X"0BFFF555FFDB9B0154150C008000E05500A4E900607F808E0000000000000000"
    , INIT_01   => X"F4FFFFF556230057A8005CAAEF150055FFFFF775C1C010E818FC4F00FEFF3900"
    , INIT_02   => X"3F0A000000005C00807FF0575040FDF759FFAB1CA2E1FCFF3F087FE5FFFF1F00"
    , INIT_03   => X"25000000F0DA03405515550700D0007B3F0000FEFCB2FC011F80783E9F00020F"
    , INIT_04   => X"000080809501E0FFFF5F5F9EF4F8FF0500000020F56000E00E00D0FAAB35F003"
    , INIT_05   => X"000080A02D001CF48F178040417F00000000000000BFE2FFF17FF501E0C33F00"
    , INIT_06   => X"00002400FAB9EA3F0F17F4557F0000000000000008BFFC22F107781FBE070012"
    , INIT_07   => X"00000054A4F603E5FFF7F3FF0700000000000000003F1FE001803BF0037EE007"
    , INIT_08   => X"27FFEAABFEB76801AA2A0C000000F8A280D0FD0060FF009D1C0000F8FFFF0300"
    , INIT_09   => X"AA7FCB2AA902002B540018F0FB0A803AFFFFF634870718D020FC1F0500000000"
    , INIT_0A   => X"6F1500000000AF00F00FFA2BA8947E37AAFE57189070F8FFFFE17FE2FFFF7F00"
    , INIT_0B   => X"0200410078BD3F80AA8A2A0700A9003F0B0000FCF864F8011EC0783E1EFC0409"
    , INIT_0C   => X"000000801BFFFF3AAFAC0A0AE8E05F0000000044AA05FCFF070078FF5FE9FF01"
    , INIT_0D   => X"000012C03B0070EA873F80AA809F000000000000007FF9FFE1FFEB01E0F1FF00"
    , INIT_0E   => X"00005001FCC7FD1F38AB8AABFF18000000000000007F8905E10F481E9E040010"
    , INIT_0F   => X"000080DA48170F2A3C3DC01C0100000000000000401F0FE0FFFF1FE001FCFF03"
    , INIT_10   => X"0AFFD5573D2710015D550E0800005C5101E4FB18007F809EE00000F0FFFF0700"
    , INIT_11   => X"F5FF949688008017BA00387E5D01505D7FFCEFB80F030CE041F81F00F0FF7F0E"
    , INIT_12   => X"9F02800000C01500FF00DD155440FFCB05FFAFB140F0F8FFFFF37FF0FFFFFF00"
    , INIT_13   => X"09000200ECC6FF4F57C515060054005F050000F8FC48A80310A0481F3EFC0108"
    , INIT_14   => X"0000008077AB00F456560102D0C02F0000000000500BF8FF0300F8FFFF57FD00"
    , INIT_15   => X"000060842F00C0F583FD4055400F00000000000000B7FCFFE1FFF703F0F9FF01"
    , INIT_16   => X"0000000AF83DFF0FE05781FE3F2100000000000020FF1003A10A402211040010"
    , INIT_17   => X"8ED900B0A8177850F1FA7FEC0000000000000008802F0FE0FFFF0FE001F8FF01"
    , INIT_18   => X"17FFABBFDA080280ABEA0721C0002F2082D0FBE1007E413D8C07000000000000"
    , INIT_19   => X"EA3F29290100C00B7D00B8AF2F00A92EBFF1FF90170C04D085F03F00E0FFFF1C"
    , INIT_1A   => X"2F05000400F002F00FA0E20BBAA47E0383364F6A076CF0FFFFFF7FF0FFFFFF01"
    , INIT_1B   => X"02000000C2030EFFBFEA0A1C00E9002D0B0000F05A9050031254401F3CFC010A"
    , INIT_1C   => X"00000080FF070AE82BAA0013A0800500000000002256F8FF0100F801E0FF7F00"
    , INIT_1D   => X"0000C4483F0080FB83CA472AA017000000000000005FFEFFC1FFEF03F0FCFF03"
    , INIT_1E   => X"00000211F5EBF82B80AF00FE4F00000000000000407F21264115402088060014"
    , INIT_1F   => X"50AA00A8502FE0A3AAFFDF5F0000000000000020001F4FE5FFFF07C000F0FF00"
    , INIT_20   => X"8BFF577DED21045155800B8444C3175041E8FF0001B8413A141F00E0FFFFCF00"
    , INIT_21   => X"FD4FCA280000C015BE00F0D38540D41F5FC08FC057000EA085C13F0000000000"
    , INIT_22   => X"17010049007E01FF0054D0157C50BF0305CB9C555E5A00F0C3FF78F80700F003"
    , INIT_23   => X"01000800C1011CC0FF7F15F203D4801F010000A9542000001280D00F7CFC030D"
    , INIT_24   => X"000000C0DF1C505057570022410001000000000008ABF07F0000F801E0F71F00"
    , INIT_25   => X"000088907F00A8FED5157F00C00D000000000000003F3EE00180DF07F87EE007"
    , INIT_26   => X"00004004EA5FE757557F01FD3F0800000000000000BF585D090048840A05001A"
    , INIT_27   => X"D0AB40E0A02B405F5595FF2F0000000000000040002FAFE2FFFF01C000C03F00"
    , INIT_28   => X"27FFAFEA0A4420A80A250E50E1FF0228ABF41E0E08C0627400FF00C0FFFF9F01"
    , INIT_29   => X"FFD490420000E0025F00FEE81290FA2F2F8007A15B0007C00903BC0700000000"
    , INIT_2A   => X"4F0000820013E00FAA0AA80BBEA57F01820031EBB03700C0073F78F80700C007"
    , INIT_2B   => X"00001080E90070A0ABFFFFBE1FAA802F00000050D80100001520E808483C800A"
    , INIT_2C   => X"000010905F70A0AABE2B00318281000000000000405F01000000000000000000"
    , INIT_2D   => X"00006240FF0055FDAAFFCC00A853000000000000005F1FE00100BE07781F800F"
    , INIT_2E   => X"00008409D4E37FBE2AF60AFD7F00000000000000207FBCAA11405450850A0015"
    , INIT_2F   => X"4EAA10E9502F80FA007AFC450000000000000040081B40050000000000000000"
    , INIT_30   => X"0AFF5F541500005D25000CAA7A7F0154D5EA053B1860237A00FE030000000000"
    , INIT_31   => X"7EA31100000070052AC07F750540F51F1700674769810BA02907801F00000000"
    , INIT_32   => X"05000005802FFE557F15D4077DD0FE01410040DFC12D00800F1E78FC0F008007"
    , INIT_33   => X"00008080C700E0415751E913FDF4801701000090B00200001A00D0F887200005"
    , INIT_34   => X"000040A05DC001F57F15001D410003000000000080BFAAAA0000000000000000"
    , INIT_35   => X"0000C4909EAAFFFFFFFFBF07D401000000000000003FBFE2A10ABC0F7C0F000F"
    , INIT_36   => X"00000812A027FEFF019C57FF9F00000000000000003F5E55A92A68A8060D000A"
    , INIT_37   => X"00000058A07F00D407A0E30A0000000000000004002FA0020000080000000000"
    , INIT_38   => X"57FF2BA2000000AE00001C55BDAA003AEBF4566D5080317400FE0700FFFF1C00"
    , INIT_39   => X"FF0702000000B80215F8F3BE0094FEAFA900D28EACC10100000E000F00000000"
    , INIT_3A   => X"92000002E0FFFFFFAB0AAA037EA57F01000080BF035900000F0C787C0F55810F"
    , INIT_3B   => X"00000080EB0080A7ABFFFF0FFAEBC00B00000080680C00800D006854D520C007"
    , INIT_3C   => X"000080D42B0007AAEF0B40818281040000000000006F05000000000000000000"
    , INIT_3D   => X"0000B0201DFFFFFF832BC8AEFA02000000000000007F7EE501107C0FBC0F001F"
    , INIT_3E   => X"0000480050FFE1FF1F78AEFD2B00000000000000005FFFFF511536F0031F800D"
    , INIT_3F   => X"00000042D08F01A83CFE7F010000000000000009545755555555250000000000"
  )
  port map (
      DI    => "00000000"
    , DIP   => "0"
    , DO    => do(2)
    , ADDR  => addr(10 downto 0)
    , CLK   => clk
    , EN    => en(2)
    , WE    => '0'
    , SSR   => '0'
  );

  ram3 : RAMB16_S9
  generic map (
      write_mode => "READ_FIRST"      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    , INIT_00   => X"0808080B0B0B08080808084828284848282948480D2818080808080101010101"
    , INIT_01   => X"08080819191908080808393928283828680D2838282848080B0B0B1919010101"
    , INIT_02   => X"080B19193B1908080839392F292817172829161528282808080B0B1919010101"
    , INIT_03   => X"08080B0B191968686828292929281017393A3A10280B2801080B191919010101"
    , INIT_04   => X"0808080808084D29292828484828483869393338280D29010801010101010101"
    , INIT_05   => X"08080808080848080829284848080839282829100F0D29594101010101010000"
    , INIT_06   => X"0808080808081008682838383A69292928182828070D08484141010100000000"
    , INIT_07   => X"080808080B083818682838381069292929182828070508484141010101010101"
    , INIT_08   => X"0808080808083838683828383A2A28292903080707054D480101010101010101"
    , INIT_09   => X"0808080808080838383A323A323202291928680541054D480505010D0D010101"
    , INIT_0A   => X"08080828686868682931303832021029192868054105454D0D0D0D0D0D0D0101"
    , INIT_0B   => X"0838382828286868290E303032101029194848284105050D48410D0541414101"
    , INIT_0C   => X"6868686969294868292930301010102919483838054505054848410141414101"
    , INIT_0D   => X"08012929292948282929383832321031194838070505050D0848020101010101"
    , INIT_0E   => X"0829292929294810152A383832323228383039050505050D0501020201010101"
    , INIT_0F   => X"080D290D2828103832323A3A323A3A393A3239050505050F0501010505050505"
    , INIT_10   => X"082929292838383232323032323830323E322905050705070D05050505050505"
    , INIT_11   => X"01293D3D3D3D3A3237323A32323232320E0A290F0F0707070D0D0D0505050505"
    , INIT_12   => X"29393D3D3B3B3A3A323232323732320A6179794D0D0F47474747474747474747"
    , INIT_13   => X"39383D393B383A3232323230383210617C78797D690D45454505454545454545"
    , INIT_14   => X"383D3D393B3A3A3232323A3B58027A787878797D7D4F0E060606060606060606"
    , INIT_15   => X"383D3D29383832323A32385958787D787878797D7D4F47474747474747474747"
    , INIT_16   => X"383D3D2F2830323A3A323218787D78787878797D7D4F45454545454545454545"
    , INIT_17   => X"38383D3D2938323232323278787D78787879797D7D4F06060606060606060606"
  )
  port map (
      DI    => "00000000"
    , DIP   => "0"
    , DO    => do(3)
    , ADDR  => addr(10 downto 0)
    , CLK   => clk
    , EN    => en(3)
    , WE    => '0'
    , SSR   => '0'
  );

end Behavioral;
